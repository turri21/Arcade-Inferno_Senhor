library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity inferno_bank_d is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of inferno_bank_d is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"0F",X"05",X"59",X"05",X"65",X"05",X"71",X"05",X"7D",X"05",X"89",X"05",X"95",
		X"05",X"A1",X"04",X"ED",X"04",X"F9",X"05",X"05",X"05",X"11",X"05",X"1D",X"05",X"29",X"05",X"35",
		X"04",X"81",X"04",X"8D",X"04",X"99",X"04",X"A5",X"04",X"B1",X"04",X"BD",X"04",X"C9",X"04",X"15",
		X"04",X"21",X"04",X"2D",X"04",X"39",X"04",X"45",X"04",X"51",X"04",X"5D",X"0C",X"01",X"0C",X"0D",
		X"0C",X"19",X"00",X"0F",X"07",X"09",X"07",X"15",X"07",X"21",X"07",X"2D",X"07",X"39",X"07",X"45",
		X"07",X"51",X"06",X"9D",X"06",X"A9",X"06",X"B5",X"06",X"C1",X"06",X"CD",X"06",X"D9",X"06",X"E5",
		X"06",X"31",X"06",X"3D",X"06",X"49",X"06",X"55",X"06",X"61",X"06",X"6D",X"06",X"79",X"05",X"C5",
		X"05",X"D1",X"05",X"DD",X"05",X"E9",X"05",X"F5",X"06",X"01",X"06",X"0D",X"0C",X"25",X"0C",X"31",
		X"0C",X"3D",X"00",X"0F",X"0E",X"71",X"0E",X"7D",X"0E",X"89",X"0E",X"95",X"0E",X"A1",X"0E",X"AD",
		X"0E",X"B9",X"0E",X"05",X"0E",X"11",X"0E",X"1D",X"0E",X"29",X"0E",X"35",X"0E",X"41",X"0E",X"4D",
		X"0D",X"81",X"0D",X"8D",X"0D",X"99",X"0D",X"A5",X"0D",X"B1",X"0D",X"BD",X"0D",X"C9",X"0D",X"15",
		X"0D",X"21",X"0D",X"2D",X"0D",X"39",X"0D",X"45",X"0D",X"51",X"0D",X"5D",X"0D",X"ED",X"0D",X"F9",
		X"00",X"0F",X"0F",X"55",X"0F",X"61",X"0F",X"6D",X"0F",X"79",X"0F",X"85",X"0F",X"91",X"0F",X"9D",
		X"10",X"15",X"10",X"21",X"10",X"2D",X"10",X"39",X"10",X"45",X"10",X"51",X"10",X"5D",X"0E",X"F5",
		X"0F",X"01",X"0F",X"0D",X"0F",X"19",X"0F",X"25",X"0F",X"31",X"0F",X"3D",X"0F",X"B5",X"0F",X"C1",
		X"0F",X"CD",X"0F",X"D9",X"0F",X"E5",X"0F",X"F1",X"0F",X"FD",X"0E",X"DD",X"0E",X"E9",X"00",X"0F",
		X"10",X"ED",X"10",X"F9",X"11",X"05",X"11",X"11",X"11",X"1D",X"11",X"29",X"11",X"35",X"11",X"AD",
		X"11",X"B9",X"11",X"C5",X"11",X"D1",X"11",X"DD",X"11",X"E9",X"11",X"F5",X"10",X"8D",X"10",X"99",
		X"10",X"A5",X"10",X"B1",X"10",X"BD",X"10",X"C9",X"10",X"D5",X"11",X"4D",X"11",X"59",X"11",X"65",
		X"11",X"71",X"11",X"7D",X"11",X"89",X"11",X"95",X"10",X"75",X"10",X"81",X"05",X"AD",X"05",X"41",
		X"04",X"D5",X"04",X"69",X"05",X"B9",X"05",X"4D",X"04",X"E1",X"04",X"75",X"07",X"5D",X"06",X"F1",
		X"06",X"85",X"06",X"19",X"07",X"69",X"06",X"FD",X"06",X"91",X"06",X"25",X"0E",X"C5",X"0E",X"59",
		X"0D",X"D5",X"0D",X"69",X"0E",X"D1",X"0E",X"65",X"0D",X"E1",X"0D",X"75",X"0F",X"A9",X"10",X"69",
		X"0F",X"49",X"10",X"09",X"0E",X"D1",X"0E",X"65",X"0D",X"E1",X"0D",X"75",X"11",X"41",X"12",X"01",
		X"10",X"E1",X"11",X"A1",X"0E",X"D1",X"0E",X"65",X"0D",X"E1",X"0D",X"75",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"25",X"12",X"31",
		X"12",X"3D",X"12",X"49",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"25",X"12",X"31",
		X"12",X"3D",X"12",X"49",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"75",X"01",X"01",X"07",X"EA",X"FE",X"FF",X"07",X"EA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"9C",X"FF",X"01",X"07",X"C3",X"00",X"FF",X"07",X"C3",X"00",X"00",X"07",X"F7",X"00",X"07",
		X"00",X"00",X"00",X"00",X"07",X"8F",X"02",X"03",X"07",X"9C",X"00",X"00",X"07",X"D0",X"00",X"07",
		X"00",X"00",X"00",X"00",X"07",X"B6",X"FE",X"03",X"07",X"75",X"00",X"00",X"07",X"82",X"00",X"08",
		X"08",X"04",X"FE",X"0D",X"00",X"00",X"00",X"00",X"07",X"EA",X"FF",X"F6",X"07",X"A9",X"00",X"08",
		X"07",X"DD",X"01",X"0D",X"00",X"00",X"00",X"00",X"07",X"C3",X"FF",X"F6",X"0C",X"CD",X"0C",X"D9",
		X"0C",X"E5",X"0C",X"F1",X"0C",X"FD",X"0D",X"09",X"0C",X"85",X"0C",X"91",X"0C",X"9D",X"0C",X"A9",
		X"0C",X"B5",X"0C",X"C1",X"00",X"0F",X"08",X"F5",X"08",X"E9",X"08",X"DD",X"08",X"D1",X"08",X"C5",
		X"08",X"B9",X"08",X"AD",X"08",X"A1",X"08",X"95",X"08",X"89",X"08",X"1D",X"09",X"01",X"00",X"00",
		X"0A",X"45",X"0A",X"15",X"09",X"55",X"09",X"25",X"0A",X"51",X"0A",X"5D",X"0A",X"69",X"0A",X"21",
		X"0A",X"2D",X"0A",X"39",X"09",X"61",X"09",X"6D",X"09",X"79",X"09",X"31",X"09",X"3D",X"09",X"49",
		X"09",X"E5",X"09",X"F1",X"09",X"FD",X"0A",X"09",X"09",X"0D",X"09",X"0D",X"09",X"B5",X"09",X"C1",
		X"09",X"CD",X"09",X"D9",X"09",X"85",X"09",X"91",X"09",X"9D",X"09",X"A9",X"08",X"59",X"08",X"65",
		X"08",X"71",X"08",X"7D",X"08",X"29",X"08",X"35",X"08",X"41",X"08",X"4D",X"00",X"0F",X"0B",X"DD",
		X"0B",X"B9",X"0B",X"05",X"0A",X"E1",X"0B",X"E9",X"0B",X"C5",X"0B",X"11",X"0A",X"ED",X"0B",X"35",
		X"0B",X"29",X"0B",X"35",X"0B",X"29",X"0A",X"B1",X"0A",X"BD",X"0A",X"C9",X"0A",X"D5",X"0B",X"95",
		X"0B",X"A1",X"0B",X"AD",X"0A",X"A5",X"0A",X"75",X"0A",X"81",X"0A",X"8D",X"0A",X"99",X"0B",X"89",
		X"0B",X"4D",X"0B",X"59",X"0B",X"65",X"0B",X"71",X"0B",X"7D",X"0B",X"41",X"0B",X"4D",X"0B",X"59",
		X"0B",X"65",X"0B",X"71",X"0B",X"7D",X"0C",X"49",X"0C",X"55",X"0C",X"61",X"0C",X"6D",X"0C",X"79",
		X"00",X"0F",X"03",X"FD",X"04",X"09",X"03",X"E5",X"03",X"F1",X"03",X"CD",X"03",X"D9",X"03",X"85",
		X"03",X"91",X"03",X"9D",X"03",X"A9",X"03",X"B5",X"03",X"C1",X"03",X"55",X"03",X"61",X"03",X"6D",
		X"03",X"79",X"08",X"11",X"12",X"0D",X"12",X"19",X"20",X"49",X"4E",X"46",X"45",X"52",X"4E",X"4F",
		X"20",X"2D",X"20",X"28",X"43",X"29",X"31",X"39",X"38",X"34",X"20",X"57",X"49",X"4C",X"4C",X"49",
		X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",
		X"49",X"4E",X"43",X"2E",X"20",X"02",X"27",X"00",X"37",X"00",X"00",X"06",X"1D",X"07",X"1D",X"01",
		X"00",X"03",X"21",X"00",X"E5",X"00",X"00",X"0A",X"17",X"0A",X"17",X"00",X"00",X"03",X"21",X"01",
		X"CB",X"00",X"00",X"08",X"17",X"08",X"17",X"00",X"00",X"04",X"27",X"02",X"83",X"00",X"00",X"07",
		X"1C",X"07",X"1C",X"00",X"00",X"05",X"21",X"03",X"47",X"00",X"00",X"0C",X"0E",X"0C",X"0E",X"00",
		X"00",X"04",X"21",X"03",X"EF",X"00",X"00",X"0C",X"11",X"0C",X"11",X"00",X"00",X"03",X"27",X"04",
		X"BB",X"00",X"00",X"06",X"1D",X"06",X"1D",X"00",X"00",X"06",X"21",X"05",X"69",X"00",X"00",X"0A",
		X"17",X"0A",X"17",X"00",X"00",X"04",X"21",X"06",X"4F",X"00",X"00",X"08",X"17",X"08",X"17",X"00",
		X"00",X"02",X"27",X"07",X"07",X"00",X"00",X"07",X"1C",X"08",X"1C",X"01",X"00",X"06",X"21",X"07",
		X"CB",X"00",X"00",X"0C",X"0E",X"0C",X"0E",X"00",X"00",X"07",X"21",X"08",X"73",X"00",X"00",X"0C",
		X"11",X"0C",X"11",X"00",X"00",X"09",X"21",X"09",X"3F",X"00",X"00",X"11",X"0E",X"11",X"0E",X"00",
		X"00",X"04",X"21",X"0A",X"2D",X"00",X"00",X"0C",X"11",X"0C",X"11",X"00",X"00",X"07",X"21",X"0A",
		X"F9",X"00",X"00",X"11",X"0E",X"11",X"0E",X"00",X"00",X"07",X"21",X"0B",X"E7",X"00",X"00",X"0C",
		X"11",X"0C",X"11",X"00",X"00",X"03",X"19",X"0C",X"B3",X"00",X"00",X"07",X"0D",X"0A",X"1D",X"02",
		X"10",X"02",X"19",X"0D",X"0E",X"00",X"00",X"06",X"0C",X"0A",X"1C",X"03",X"10",X"02",X"18",X"0D",
		X"56",X"00",X"00",X"06",X"0D",X"0A",X"1E",X"03",X"11",X"03",X"18",X"0D",X"A4",X"00",X"00",X"07",
		X"0C",X"0A",X"1D",X"02",X"11",X"04",X"18",X"0D",X"F8",X"00",X"00",X"08",X"0C",X"0A",X"1D",X"01",
		X"11",X"02",X"18",X"0E",X"58",X"00",X"00",X"07",X"0C",X"0A",X"1D",X"03",X"11",X"02",X"18",X"0E",
		X"AC",X"00",X"00",X"05",X"0C",X"0A",X"1D",X"03",X"11",X"03",X"22",X"0E",X"E8",X"00",X"00",X"07",
		X"0B",X"0A",X"12",X"02",X"07",X"02",X"29",X"0F",X"35",X"00",X"00",X"07",X"12",X"0A",X"12",X"03",
		X"00",X"03",X"19",X"0F",X"B3",X"00",X"00",X"07",X"0D",X"0A",X"1D",X"02",X"10",X"03",X"19",X"10",
		X"0E",X"00",X"00",X"06",X"0C",X"0A",X"1C",X"02",X"10",X"03",X"18",X"10",X"56",X"00",X"00",X"06",
		X"0D",X"0A",X"1E",X"02",X"11",X"03",X"18",X"10",X"A4",X"00",X"00",X"07",X"0C",X"0A",X"1D",X"02",
		X"11",X"03",X"18",X"10",X"F8",X"00",X"00",X"08",X"0C",X"0A",X"1D",X"02",X"11",X"04",X"18",X"11",
		X"58",X"00",X"00",X"07",X"0C",X"0A",X"1D",X"01",X"11",X"02",X"18",X"11",X"AC",X"00",X"00",X"05",
		X"0C",X"0A",X"1D",X"03",X"11",X"03",X"22",X"11",X"E8",X"00",X"00",X"07",X"0B",X"0A",X"12",X"02",
		X"07",X"04",X"29",X"12",X"35",X"00",X"00",X"07",X"12",X"0A",X"12",X"01",X"00",X"02",X"17",X"12",
		X"B3",X"00",X"00",X"05",X"0D",X"0A",X"1F",X"03",X"12",X"03",X"18",X"12",X"F4",X"00",X"00",X"06",
		X"0D",X"0A",X"1E",X"02",X"11",X"04",X"17",X"13",X"42",X"00",X"00",X"09",X"0C",X"0A",X"1E",X"01",
		X"12",X"02",X"17",X"13",X"AE",X"00",X"00",X"05",X"0C",X"0A",X"1E",X"03",X"12",X"03",X"18",X"13",
		X"EA",X"00",X"00",X"05",X"0F",X"0A",X"20",X"02",X"11",X"03",X"17",X"14",X"35",X"00",X"00",X"06",
		X"0E",X"0A",X"20",X"02",X"12",X"02",X"17",X"14",X"89",X"00",X"00",X"05",X"0D",X"0A",X"1F",X"03",
		X"12",X"03",X"22",X"14",X"CA",X"00",X"00",X"07",X"0B",X"0A",X"12",X"02",X"07",X"03",X"29",X"15",
		X"17",X"00",X"00",X"07",X"12",X"0A",X"12",X"02",X"00",X"02",X"17",X"15",X"95",X"00",X"00",X"05",
		X"0D",X"0A",X"1F",X"03",X"12",X"02",X"18",X"15",X"D6",X"00",X"00",X"06",X"0D",X"0A",X"1E",X"03",
		X"11",X"04",X"17",X"16",X"24",X"00",X"00",X"09",X"0C",X"0A",X"1E",X"01",X"12",X"02",X"17",X"16",
		X"90",X"00",X"00",X"05",X"0C",X"0A",X"1E",X"03",X"12",X"01",X"18",X"16",X"CC",X"00",X"00",X"05",
		X"0F",X"0A",X"20",X"04",X"11",X"02",X"17",X"17",X"17",X"00",X"00",X"06",X"0E",X"0A",X"20",X"03",
		X"12",X"02",X"17",X"17",X"6B",X"00",X"00",X"05",X"0D",X"0A",X"1F",X"03",X"12",X"03",X"22",X"17",
		X"AC",X"00",X"00",X"07",X"0B",X"0A",X"12",X"02",X"07",X"03",X"29",X"17",X"F9",X"00",X"00",X"07",
		X"12",X"0A",X"12",X"02",X"00",X"03",X"19",X"18",X"77",X"00",X"00",X"07",X"0E",X"0A",X"1B",X"02",
		X"0D",X"02",X"19",X"18",X"D9",X"00",X"00",X"06",X"0C",X"0A",X"19",X"03",X"0D",X"02",X"18",X"19",
		X"21",X"00",X"00",X"06",X"0D",X"0A",X"1B",X"03",X"0E",X"03",X"18",X"19",X"6F",X"00",X"00",X"07",
		X"0C",X"0A",X"1A",X"02",X"0E",X"04",X"18",X"19",X"C3",X"00",X"00",X"08",X"0C",X"0A",X"1A",X"01",
		X"0E",X"02",X"18",X"1A",X"23",X"00",X"00",X"07",X"0C",X"0A",X"1A",X"03",X"0E",X"02",X"18",X"1A",
		X"77",X"00",X"00",X"05",X"0C",X"0A",X"1A",X"03",X"0E",X"04",X"22",X"1A",X"B3",X"00",X"00",X"08",
		X"0B",X"0A",X"0F",X"01",X"04",X"04",X"26",X"1B",X"0B",X"00",X"00",X"07",X"0F",X"0A",X"0F",X"01",
		X"00",X"03",X"19",X"1B",X"74",X"00",X"00",X"07",X"0E",X"0A",X"1B",X"02",X"0D",X"03",X"19",X"1B",
		X"D6",X"00",X"00",X"06",X"0C",X"0A",X"19",X"02",X"0D",X"03",X"18",X"1C",X"1E",X"00",X"00",X"06",
		X"0D",X"0A",X"1B",X"02",X"0E",X"03",X"18",X"1C",X"6C",X"00",X"00",X"07",X"0C",X"0A",X"1A",X"02",
		X"0E",X"03",X"18",X"1C",X"C0",X"00",X"00",X"08",X"0C",X"0A",X"1A",X"02",X"0E",X"04",X"18",X"1D",
		X"20",X"00",X"00",X"07",X"0C",X"0A",X"1A",X"01",X"0E",X"02",X"18",X"1D",X"74",X"00",X"00",X"05",
		X"0C",X"0A",X"1A",X"03",X"0E",X"03",X"22",X"1D",X"B0",X"00",X"00",X"08",X"0B",X"0A",X"0F",X"02",
		X"04",X"02",X"26",X"1E",X"08",X"00",X"00",X"07",X"0F",X"0A",X"0F",X"03",X"00",X"02",X"17",X"1E",
		X"71",X"00",X"00",X"05",X"0D",X"0A",X"1C",X"03",X"0F",X"03",X"18",X"1E",X"B2",X"00",X"00",X"06",
		X"0D",X"0A",X"1B",X"02",X"0E",X"04",X"17",X"1F",X"00",X"00",X"00",X"09",X"0C",X"0A",X"1B",X"01",
		X"0F",X"02",X"17",X"1F",X"6C",X"00",X"00",X"05",X"0C",X"0A",X"1B",X"03",X"0F",X"03",X"18",X"1F",
		X"A8",X"00",X"00",X"05",X"0F",X"0A",X"1D",X"02",X"0E",X"03",X"17",X"1F",X"F3",X"00",X"00",X"06",
		X"0E",X"0A",X"1D",X"02",X"0F",X"02",X"17",X"20",X"47",X"00",X"00",X"05",X"0D",X"0A",X"1C",X"03",
		X"0F",X"03",X"22",X"20",X"88",X"00",X"00",X"07",X"0B",X"0A",X"0F",X"02",X"04",X"03",X"26",X"20",
		X"D5",X"00",X"00",X"07",X"0F",X"0A",X"0F",X"02",X"00",X"02",X"17",X"21",X"3E",X"00",X"00",X"05",
		X"0D",X"0A",X"1C",X"03",X"0F",X"02",X"18",X"21",X"7F",X"00",X"00",X"06",X"0D",X"0A",X"1B",X"03",
		X"0E",X"04",X"17",X"21",X"CD",X"00",X"00",X"09",X"0C",X"0A",X"1B",X"01",X"0F",X"02",X"17",X"22",
		X"39",X"00",X"00",X"05",X"0C",X"0A",X"1B",X"03",X"0F",X"01",X"18",X"22",X"75",X"00",X"00",X"05",
		X"0F",X"0A",X"1D",X"04",X"0E",X"02",X"17",X"22",X"C0",X"00",X"00",X"06",X"0E",X"0A",X"1D",X"03",
		X"0F",X"02",X"17",X"23",X"14",X"00",X"00",X"05",X"0D",X"0A",X"1C",X"03",X"0F",X"03",X"22",X"23",
		X"55",X"00",X"00",X"07",X"0B",X"0A",X"0F",X"02",X"04",X"03",X"26",X"23",X"A2",X"00",X"00",X"07",
		X"0F",X"0A",X"0F",X"02",X"00",X"03",X"0E",X"7A",X"34",X"FD",X"04",X"04",X"04",X"07",X"82",X"07",
		X"8F",X"00",X"03",X"0D",X"7A",X"44",X"FD",X"04",X"03",X"07",X"07",X"8F",X"07",X"8F",X"F8",X"05",
		X"07",X"7A",X"59",X"FD",X"04",X"03",X"06",X"07",X"8F",X"07",X"8F",X"F8",X"00",X"0E",X"7A",X"6B",
		X"03",X"04",X"04",X"04",X"07",X"A9",X"07",X"B6",X"00",X"FF",X"0D",X"7A",X"7B",X"03",X"04",X"03",
		X"07",X"07",X"B6",X"07",X"B6",X"F8",X"FD",X"07",X"7A",X"90",X"03",X"04",X"03",X"06",X"07",X"B6",
		X"07",X"B6",X"F8",X"03",X"13",X"7A",X"A2",X"FC",X"FC",X"04",X"04",X"07",X"D0",X"07",X"DD",X"00",
		X"03",X"16",X"7A",X"B2",X"FC",X"FC",X"03",X"06",X"07",X"DD",X"07",X"DD",X"F8",X"05",X"1C",X"7A",
		X"C4",X"FC",X"FC",X"03",X"06",X"07",X"DD",X"07",X"DD",X"F8",X"00",X"13",X"7A",X"D6",X"02",X"FC",
		X"04",X"04",X"07",X"F7",X"08",X"04",X"00",X"FF",X"16",X"7A",X"E6",X"02",X"FC",X"03",X"06",X"08",
		X"04",X"08",X"04",X"F8",X"FD",X"1C",X"7A",X"F8",X"02",X"FC",X"03",X"06",X"08",X"04",X"08",X"04",
		X"F8",X"02",X"11",X"24",X"0B",X"00",X"00",X"05",X"05",X"0A",X"1D",X"03",X"18",X"05",X"17",X"24",
		X"24",X"00",X"1B",X"0B",X"0D",X"0C",X"19",X"01",X"0C",X"03",X"16",X"24",X"B3",X"00",X"1B",X"06",
		X"07",X"0C",X"14",X"03",X"0D",X"05",X"19",X"24",X"DD",X"00",X"1B",X"09",X"0D",X"0C",X"17",X"01",
		X"0A",X"06",X"1A",X"25",X"52",X"00",X"1B",X"0C",X"0F",X"0C",X"18",X"00",X"09",X"06",X"1A",X"26",
		X"06",X"00",X"1B",X"0C",X"11",X"0C",X"1A",X"00",X"09",X"03",X"16",X"26",X"D2",X"00",X"1B",X"06",
		X"07",X"0C",X"14",X"03",X"0D",X"04",X"19",X"26",X"FC",X"00",X"1B",X"09",X"0D",X"0C",X"17",X"02",
		X"0A",X"06",X"1A",X"27",X"71",X"00",X"1B",X"0C",X"0F",X"0C",X"18",X"00",X"09",X"06",X"1A",X"28",
		X"25",X"00",X"1B",X"0C",X"11",X"0C",X"1A",X"00",X"09",X"06",X"1A",X"28",X"F1",X"00",X"1B",X"0C",
		X"11",X"0C",X"1A",X"00",X"09",X"06",X"1A",X"29",X"BD",X"00",X"1B",X"0C",X"11",X"0C",X"1A",X"00",
		X"09",X"06",X"1A",X"2A",X"C0",X"00",X"1B",X"0C",X"11",X"0C",X"1A",X"00",X"09",X"06",X"1A",X"2B",
		X"8C",X"00",X"1B",X"0C",X"11",X"0C",X"1A",X"00",X"09",X"06",X"17",X"2C",X"58",X"00",X"1B",X"0B",
		X"0F",X"0C",X"1B",X"00",X"0C",X"06",X"1A",X"2C",X"FD",X"00",X"1B",X"0C",X"11",X"0C",X"1A",X"00",
		X"09",X"06",X"1A",X"2D",X"C9",X"00",X"1B",X"0C",X"11",X"0C",X"1A",X"00",X"09",X"06",X"1A",X"2E",
		X"95",X"00",X"1B",X"0C",X"11",X"0C",X"1A",X"00",X"09",X"06",X"1A",X"2F",X"61",X"00",X"1B",X"0C",
		X"11",X"0C",X"1A",X"00",X"09",X"05",X"17",X"30",X"2D",X"00",X"1B",X"0B",X"0F",X"0C",X"1B",X"01",
		X"0C",X"03",X"1C",X"30",X"D2",X"00",X"1B",X"06",X"13",X"0C",X"1A",X"03",X"07",X"02",X"1E",X"31",
		X"44",X"00",X"1B",X"04",X"03",X"0C",X"08",X"04",X"05",X"02",X"1E",X"31",X"50",X"00",X"1B",X"04",
		X"03",X"0C",X"08",X"04",X"05",X"05",X"23",X"31",X"5C",X"00",X"1B",X"0B",X"11",X"0C",X"11",X"01",
		X"00",X"08",X"16",X"32",X"17",X"00",X"1B",X"05",X"04",X"0E",X"11",X"00",X"0D",X"0A",X"16",X"32",
		X"2B",X"00",X"1B",X"07",X"07",X"10",X"14",X"00",X"0D",X"0B",X"17",X"32",X"5C",X"00",X"1B",X"08",
		X"09",X"11",X"15",X"00",X"0C",X"06",X"23",X"32",X"A4",X"00",X"1B",X"0B",X"11",X"0C",X"11",X"00",
		X"00",X"FD",X"16",X"33",X"5F",X"00",X"1B",X"05",X"04",X"0E",X"11",X"09",X"0D",X"FD",X"16",X"33",
		X"73",X"00",X"1B",X"07",X"07",X"10",X"14",X"09",X"0D",X"FD",X"17",X"33",X"A4",X"00",X"1B",X"08",
		X"09",X"11",X"15",X"09",X"0C",X"05",X"25",X"33",X"EC",X"00",X"1B",X"0C",X"0F",X"0D",X"0D",X"00",
		X"FE",X"06",X"25",X"34",X"A0",X"00",X"1B",X"0E",X"11",X"0E",X"0F",X"FF",X"FE",X"06",X"25",X"35",
		X"8E",X"00",X"1B",X"0D",X"10",X"0D",X"0E",X"FF",X"FE",X"06",X"27",X"36",X"5E",X"00",X"1B",X"0D",
		X"12",X"0D",X"0E",X"FF",X"FC",X"07",X"25",X"37",X"48",X"00",X"1B",X"0C",X"0F",X"0D",X"0D",X"FF",
		X"FE",X"08",X"25",X"37",X"FC",X"00",X"1B",X"0E",X"11",X"0E",X"0F",X"FF",X"FE",X"07",X"25",X"38",
		X"EA",X"00",X"1B",X"0D",X"10",X"0D",X"0E",X"FF",X"FE",X"07",X"27",X"39",X"BA",X"00",X"1B",X"0D",
		X"12",X"0D",X"0E",X"FF",X"FC",X"01",X"25",X"3A",X"A4",X"00",X"1B",X"02",X"08",X"0C",X"06",X"04",
		X"FE",X"01",X"25",X"3A",X"B4",X"00",X"1B",X"02",X"08",X"0C",X"06",X"04",X"FE",X"01",X"25",X"3A",
		X"C4",X"00",X"1B",X"02",X"08",X"0C",X"06",X"04",X"FE",X"01",X"25",X"3A",X"D4",X"00",X"1B",X"02",
		X"08",X"0C",X"06",X"04",X"FE",X"05",X"23",X"3A",X"E4",X"00",X"1B",X"0A",X"11",X"0C",X"11",X"01",
		X"00",X"07",X"24",X"3B",X"8E",X"00",X"1B",X"04",X"04",X"0D",X"03",X"FF",X"FF",X"09",X"26",X"3B",
		X"9E",X"00",X"1B",X"07",X"07",X"0F",X"04",X"FF",X"FD",X"0A",X"28",X"3B",X"CF",X"00",X"1B",X"07",
		X"0A",X"10",X"05",X"FF",X"FB",X"05",X"23",X"3C",X"15",X"00",X"1B",X"0A",X"11",X"0C",X"11",X"01",
		X"00",X"FD",X"24",X"3C",X"BF",X"00",X"1B",X"04",X"04",X"0D",X"03",X"08",X"FF",X"FE",X"26",X"3C",
		X"CF",X"00",X"1B",X"07",X"07",X"0F",X"04",X"07",X"FD",X"FD",X"28",X"3D",X"00",X"00",X"1B",X"07",
		X"0A",X"10",X"05",X"08",X"FB",X"01",X"15",X"3D",X"46",X"0B",X"F5",X"03",X"07",X"0B",X"19",X"04",
		X"08",X"02",X"13",X"3D",X"5B",X"0B",X"F5",X"05",X"06",X"0B",X"19",X"03",X"0A",X"03",X"14",X"3D",
		X"79",X"0B",X"F5",X"07",X"08",X"0B",X"19",X"02",X"09",X"03",X"16",X"3D",X"B1",X"0B",X"F5",X"07",
		X"0B",X"0B",X"19",X"02",X"07",X"02",X"0D",X"3D",X"FE",X"0B",X"F5",X"05",X"05",X"0B",X"19",X"03",
		X"10",X"03",X"1A",X"3E",X"17",X"0B",X"F5",X"07",X"0B",X"0B",X"19",X"02",X"03",X"05",X"1D",X"3E",
		X"64",X"0B",X"F5",X"0B",X"11",X"0B",X"19",X"00",X"00",X"06",X"1F",X"3F",X"1F",X"0B",X"F5",X"0D",
		X"15",X"0D",X"19",X"00",X"00",X"08",X"21",X"40",X"30",X"0B",X"F5",X"11",X"19",X"11",X"19",X"00",
		X"00",X"08",X"15",X"42",X"81",X"0A",X"F9",X"0A",X"0D",X"0E",X"19",X"00",X"08",X"05",X"15",X"43",
		X"03",X"0A",X"F9",X"07",X"13",X"0B",X"1B",X"00",X"08",X"04",X"12",X"43",X"88",X"0A",X"F9",X"07",
		X"09",X"0B",X"19",X"01",X"0B",X"01",X"15",X"43",X"C7",X"0B",X"1D",X"0A",X"0D",X"0E",X"19",X"04",
		X"08",X"01",X"15",X"44",X"49",X"0B",X"1D",X"07",X"13",X"0B",X"1B",X"04",X"08",X"02",X"12",X"44",
		X"CE",X"0B",X"1D",X"07",X"09",X"0B",X"19",X"03",X"0B",X"03",X"15",X"45",X"0D",X"0B",X"F5",X"05",
		X"13",X"0B",X"1B",X"02",X"08",X"01",X"15",X"45",X"6C",X"0B",X"F5",X"05",X"13",X"0B",X"1B",X"04",
		X"08",X"02",X"1A",X"45",X"CB",X"0B",X"F5",X"06",X"05",X"0B",X"19",X"03",X"03",X"02",X"1B",X"45",
		X"E9",X"0B",X"F5",X"05",X"07",X"0B",X"19",X"03",X"02",X"02",X"1B",X"46",X"0C",X"0B",X"F5",X"05",
		X"0D",X"0B",X"19",X"03",X"02",X"02",X"1D",X"46",X"4D",X"0B",X"F5",X"05",X"13",X"0B",X"19",X"03",
		X"00",X"02",X"20",X"46",X"AC",X"0B",X"F5",X"05",X"1A",X"0B",X"1A",X"03",X"00",X"03",X"1F",X"47",
		X"2E",X"0B",X"F5",X"08",X"1D",X"0B",X"1D",X"02",X"00",X"03",X"1A",X"48",X"16",X"0B",X"F5",X"06",
		X"05",X"0B",X"19",X"02",X"03",X"05",X"1D",X"48",X"34",X"0B",X"F5",X"0B",X"0D",X"0B",X"19",X"00",
		X"00",X"05",X"1C",X"48",X"C3",X"0B",X"F5",X"0B",X"0C",X"0B",X"19",X"00",X"01",X"05",X"1C",X"49",
		X"47",X"0B",X"F5",X"0B",X"0C",X"0B",X"19",X"00",X"01",X"07",X"21",X"4A",X"65",X"0B",X"D1",X"09",
		X"10",X"0D",X"19",X"00",X"00",X"07",X"16",X"4A",X"F5",X"0B",X"D1",X"09",X"0A",X"0D",X"19",X"00",
		X"07",X"04",X"14",X"4B",X"86",X"0B",X"D1",X"07",X"09",X"0B",X"19",X"01",X"09",X"01",X"21",X"4B",
		X"C5",X"0B",X"F5",X"09",X"10",X"0D",X"19",X"04",X"00",X"01",X"16",X"4C",X"55",X"0B",X"F5",X"09",
		X"0A",X"0D",X"19",X"04",X"07",X"02",X"14",X"4C",X"AF",X"0B",X"F5",X"07",X"09",X"0B",X"19",X"03",
		X"09",X"05",X"18",X"4C",X"EE",X"00",X"00",X"0B",X"13",X"0B",X"24",X"00",X"11",X"05",X"19",X"4D",
		X"BF",X"00",X"00",X"0B",X"15",X"0B",X"25",X"00",X"10",X"04",X"17",X"4E",X"A6",X"00",X"00",X"09",
		X"11",X"0A",X"23",X"01",X"12",X"05",X"18",X"4F",X"3F",X"00",X"00",X"0B",X"13",X"0B",X"21",X"00",
		X"0E",X"05",X"19",X"50",X"10",X"00",X"00",X"0B",X"15",X"0B",X"22",X"00",X"0D",X"04",X"17",X"50",
		X"F7",X"00",X"00",X"09",X"11",X"0A",X"20",X"01",X"0F",X"03",X"23",X"51",X"90",X"00",X"00",X"07",
		X"19",X"0A",X"1F",X"02",X"06",X"03",X"23",X"52",X"3F",X"00",X"00",X"07",X"19",X"0A",X"1F",X"02",
		X"06",X"03",X"23",X"52",X"EE",X"00",X"00",X"07",X"19",X"0A",X"1F",X"02",X"06",X"03",X"23",X"53",
		X"9D",X"00",X"00",X"07",X"19",X"0A",X"1F",X"02",X"06",X"03",X"13",X"54",X"4C",X"00",X"00",X"07",
		X"09",X"0A",X"1F",X"02",X"16",X"03",X"20",X"54",X"8B",X"00",X"00",X"06",X"07",X"06",X"09",X"00",
		X"02",X"03",X"20",X"54",X"B5",X"00",X"00",X"06",X"07",X"06",X"09",X"00",X"02",X"02",X"1F",X"54",
		X"DF",X"00",X"00",X"05",X"06",X"05",X"09",X"00",X"03",X"02",X"20",X"54",X"FD",X"00",X"00",X"06",
		X"07",X"06",X"09",X"00",X"02",X"02",X"20",X"55",X"27",X"00",X"00",X"06",X"07",X"06",X"09",X"00",
		X"02",X"02",X"1F",X"55",X"51",X"00",X"00",X"05",X"06",X"05",X"09",X"00",X"03",X"03",X"20",X"55",
		X"6F",X"00",X"00",X"06",X"07",X"06",X"09",X"00",X"02",X"03",X"20",X"55",X"99",X"00",X"00",X"06",
		X"07",X"06",X"09",X"00",X"02",X"02",X"20",X"55",X"C3",X"00",X"00",X"05",X"06",X"05",X"08",X"00",
		X"02",X"02",X"20",X"55",X"E1",X"00",X"00",X"06",X"07",X"06",X"09",X"00",X"02",X"02",X"20",X"56",
		X"0B",X"00",X"00",X"06",X"07",X"06",X"09",X"00",X"02",X"02",X"20",X"56",X"35",X"00",X"00",X"05",
		X"06",X"05",X"08",X"00",X"02",X"03",X"1C",X"56",X"53",X"00",X"00",X"06",X"0F",X"09",X"16",X"01",
		X"07",X"03",X"1C",X"56",X"AD",X"00",X"00",X"07",X"0E",X"09",X"15",X"01",X"07",X"02",X"1C",X"57",
		X"0F",X"00",X"00",X"06",X"11",X"09",X"18",X"02",X"07",X"03",X"1C",X"57",X"75",X"00",X"00",X"06",
		X"0F",X"09",X"16",X"01",X"07",X"03",X"1C",X"57",X"CF",X"00",X"00",X"07",X"0F",X"09",X"16",X"01",
		X"07",X"02",X"1C",X"58",X"38",X"00",X"00",X"06",X"10",X"09",X"17",X"02",X"07",X"03",X"1B",X"58",
		X"98",X"00",X"00",X"07",X"0E",X"09",X"16",X"01",X"08",X"02",X"23",X"58",X"FA",X"00",X"00",X"06",
		X"0A",X"09",X"0A",X"02",X"00",X"03",X"23",X"59",X"36",X"00",X"00",X"07",X"0A",X"09",X"0A",X"01",
		X"00",X"02",X"1C",X"59",X"7C",X"00",X"00",X"06",X"0F",X"09",X"16",X"02",X"07",X"03",X"1C",X"59",
		X"D6",X"00",X"00",X"07",X"0E",X"09",X"15",X"01",X"07",X"03",X"1C",X"5A",X"38",X"00",X"00",X"06",
		X"11",X"09",X"18",X"01",X"07",X"02",X"1C",X"5A",X"9E",X"00",X"00",X"06",X"0F",X"09",X"16",X"02",
		X"07",X"03",X"1C",X"5A",X"F8",X"00",X"00",X"07",X"0F",X"09",X"16",X"01",X"07",X"03",X"1C",X"5B",
		X"61",X"00",X"00",X"06",X"10",X"09",X"17",X"01",X"07",X"03",X"1B",X"5B",X"C1",X"00",X"00",X"07",
		X"0E",X"09",X"16",X"01",X"08",X"03",X"23",X"5C",X"23",X"00",X"00",X"06",X"0A",X"09",X"0A",X"01",
		X"00",X"03",X"23",X"5C",X"5F",X"00",X"00",X"07",X"0A",X"09",X"0A",X"01",X"00",X"01",X"1E",X"5C",
		X"A5",X"00",X"00",X"03",X"05",X"09",X"0A",X"03",X"05",X"01",X"1E",X"5C",X"B4",X"00",X"00",X"03",
		X"05",X"09",X"0A",X"03",X"05",X"02",X"1A",X"5C",X"C3",X"00",X"00",X"06",X"0F",X"09",X"18",X"02",
		X"09",X"03",X"19",X"5D",X"1D",X"00",X"00",X"06",X"0C",X"09",X"16",X"01",X"0A",X"03",X"1A",X"5D",
		X"65",X"00",X"00",X"07",X"0D",X"09",X"16",X"01",X"09",X"02",X"1A",X"5D",X"C0",X"00",X"00",X"07",
		X"0F",X"09",X"18",X"02",X"09",X"03",X"1A",X"5E",X"29",X"00",X"00",X"07",X"0E",X"09",X"17",X"01",
		X"09",X"03",X"1A",X"5E",X"8B",X"00",X"00",X"07",X"0F",X"09",X"18",X"01",X"09",X"04",X"1A",X"5E",
		X"F4",X"00",X"00",X"08",X"0E",X"09",X"17",X"00",X"09",X"02",X"23",X"5F",X"64",X"00",X"00",X"05",
		X"0A",X"09",X"0A",X"02",X"00",X"04",X"21",X"5F",X"96",X"00",X"00",X"08",X"08",X"09",X"0A",X"00",
		X"02",X"03",X"1A",X"5F",X"D6",X"00",X"00",X"06",X"0F",X"09",X"18",X"01",X"09",X"02",X"19",X"60",
		X"30",X"00",X"00",X"06",X"0C",X"09",X"16",X"02",X"0A",X"03",X"1A",X"60",X"78",X"00",X"00",X"07",
		X"0D",X"09",X"16",X"01",X"09",X"04",X"1A",X"60",X"D3",X"00",X"00",X"07",X"0F",X"09",X"18",X"00",
		X"09",X"03",X"1A",X"61",X"3C",X"00",X"00",X"07",X"0E",X"09",X"17",X"01",X"09",X"03",X"1A",X"61",
		X"9E",X"00",X"00",X"07",X"0F",X"09",X"18",X"01",X"09",X"03",X"1A",X"62",X"07",X"00",X"00",X"08",
		X"0E",X"09",X"17",X"01",X"09",X"02",X"23",X"62",X"77",X"00",X"00",X"05",X"0A",X"09",X"0A",X"02",
		X"00",X"03",X"21",X"62",X"A9",X"00",X"00",X"08",X"08",X"09",X"0A",X"01",X"02",X"01",X"1E",X"62",
		X"E9",X"00",X"00",X"03",X"05",X"09",X"0A",X"03",X"05",X"01",X"1E",X"62",X"F8",X"00",X"00",X"03",
		X"05",X"09",X"0A",X"03",X"05",X"02",X"1C",X"63",X"07",X"00",X"00",X"06",X"0F",X"09",X"16",X"02",
		X"07",X"03",X"1C",X"63",X"61",X"00",X"00",X"07",X"0E",X"09",X"15",X"01",X"07",X"03",X"1C",X"63",
		X"C3",X"00",X"00",X"06",X"11",X"09",X"18",X"01",X"07",X"02",X"1C",X"64",X"29",X"00",X"00",X"06",
		X"0F",X"09",X"16",X"02",X"07",X"03",X"1C",X"64",X"83",X"00",X"00",X"07",X"0F",X"09",X"16",X"01",
		X"07",X"03",X"1C",X"64",X"EC",X"00",X"00",X"06",X"10",X"09",X"17",X"01",X"07",X"03",X"1B",X"65",
		X"4C",X"00",X"00",X"07",X"0E",X"09",X"16",X"01",X"08",X"03",X"23",X"65",X"AE",X"00",X"00",X"06",
		X"0A",X"09",X"0A",X"01",X"00",X"03",X"1A",X"65",X"EA",X"00",X"00",X"06",X"0F",X"09",X"18",X"01",
		X"09",X"02",X"19",X"66",X"44",X"00",X"00",X"06",X"0C",X"09",X"16",X"02",X"0A",X"03",X"1A",X"66",
		X"8C",X"00",X"00",X"07",X"0D",X"09",X"16",X"01",X"09",X"04",X"1A",X"66",X"E7",X"00",X"00",X"07",
		X"0F",X"09",X"18",X"00",X"09",X"03",X"1A",X"67",X"50",X"00",X"00",X"07",X"0E",X"09",X"17",X"01",
		X"09",X"03",X"1A",X"67",X"B2",X"00",X"00",X"07",X"0F",X"09",X"18",X"01",X"09",X"03",X"1A",X"68",
		X"1B",X"00",X"00",X"08",X"0E",X"09",X"17",X"01",X"09",X"02",X"23",X"68",X"8B",X"00",X"00",X"05",
		X"0A",X"09",X"0A",X"02",X"00",X"03",X"1C",X"68",X"BD",X"00",X"00",X"06",X"0F",X"09",X"16",X"01",
		X"07",X"03",X"1C",X"69",X"17",X"00",X"00",X"07",X"0E",X"09",X"15",X"01",X"07",X"02",X"1C",X"69",
		X"79",X"00",X"00",X"06",X"11",X"09",X"18",X"02",X"07",X"03",X"1C",X"69",X"DF",X"00",X"00",X"06",
		X"0F",X"09",X"16",X"01",X"07",X"03",X"1C",X"6A",X"39",X"00",X"00",X"07",X"0F",X"09",X"16",X"01",
		X"07",X"02",X"1C",X"6A",X"A2",X"00",X"00",X"06",X"10",X"09",X"17",X"02",X"07",X"03",X"1B",X"6B",
		X"02",X"00",X"00",X"07",X"0E",X"09",X"16",X"01",X"08",X"02",X"23",X"6B",X"9B",X"00",X"00",X"06",
		X"0A",X"09",X"0A",X"02",X"00",X"02",X"1A",X"6B",X"D7",X"00",X"00",X"06",X"0F",X"09",X"18",X"02",
		X"09",X"03",X"19",X"6C",X"31",X"00",X"00",X"06",X"0C",X"09",X"16",X"01",X"0A",X"03",X"1A",X"6C",
		X"79",X"00",X"00",X"07",X"0D",X"09",X"16",X"01",X"09",X"02",X"1A",X"6C",X"D4",X"00",X"00",X"07",
		X"0F",X"09",X"18",X"02",X"09",X"03",X"1A",X"6D",X"3D",X"00",X"00",X"07",X"0E",X"09",X"17",X"01",
		X"09",X"03",X"1A",X"6D",X"9F",X"00",X"00",X"07",X"0F",X"09",X"18",X"01",X"09",X"04",X"1A",X"6E",
		X"08",X"00",X"00",X"08",X"0E",X"09",X"17",X"00",X"09",X"02",X"23",X"6E",X"78",X"00",X"00",X"05",
		X"0A",X"09",X"0A",X"02",X"00",X"01",X"1E",X"6E",X"AA",X"00",X"00",X"03",X"05",X"09",X"0A",X"03",
		X"05",X"01",X"1E",X"6E",X"B9",X"00",X"00",X"03",X"05",X"09",X"0A",X"03",X"05",X"02",X"1C",X"6E",
		X"C8",X"00",X"00",X"06",X"0F",X"09",X"16",X"02",X"07",X"03",X"1C",X"6F",X"22",X"00",X"00",X"07",
		X"0E",X"09",X"15",X"01",X"07",X"03",X"1C",X"6F",X"84",X"00",X"00",X"06",X"11",X"09",X"18",X"01",
		X"07",X"02",X"1C",X"6F",X"EA",X"00",X"00",X"06",X"0F",X"09",X"16",X"02",X"07",X"03",X"1C",X"70",
		X"44",X"00",X"00",X"07",X"0F",X"09",X"16",X"01",X"07",X"03",X"1C",X"70",X"AD",X"00",X"00",X"06",
		X"10",X"09",X"17",X"01",X"07",X"03",X"1B",X"71",X"0D",X"00",X"00",X"07",X"0E",X"09",X"16",X"01",
		X"08",X"03",X"23",X"71",X"6F",X"00",X"00",X"06",X"0A",X"09",X"0A",X"01",X"00",X"03",X"1A",X"71",
		X"AB",X"00",X"00",X"06",X"0F",X"09",X"18",X"01",X"09",X"02",X"19",X"72",X"05",X"00",X"00",X"06",
		X"0C",X"09",X"16",X"02",X"0A",X"03",X"1A",X"72",X"4D",X"00",X"00",X"07",X"0D",X"09",X"16",X"01",
		X"09",X"04",X"1A",X"72",X"A8",X"00",X"00",X"07",X"0F",X"09",X"18",X"00",X"09",X"03",X"1A",X"73",
		X"11",X"00",X"00",X"07",X"0E",X"09",X"17",X"01",X"09",X"03",X"1A",X"73",X"73",X"00",X"00",X"07",
		X"0F",X"09",X"18",X"01",X"09",X"03",X"1A",X"73",X"DC",X"00",X"00",X"08",X"0E",X"09",X"17",X"01",
		X"09",X"02",X"23",X"74",X"4C",X"00",X"00",X"05",X"0A",X"09",X"0A",X"02",X"00",X"03",X"1C",X"74",
		X"7E",X"00",X"00",X"06",X"0F",X"09",X"16",X"01",X"07",X"03",X"1C",X"74",X"D8",X"00",X"00",X"07",
		X"0E",X"09",X"15",X"01",X"07",X"02",X"1C",X"75",X"3A",X"00",X"00",X"06",X"11",X"09",X"18",X"02",
		X"07",X"03",X"1C",X"75",X"A0",X"00",X"00",X"06",X"0F",X"09",X"16",X"01",X"07",X"03",X"1C",X"75",
		X"FA",X"00",X"00",X"07",X"0F",X"09",X"16",X"01",X"07",X"02",X"1C",X"76",X"63",X"00",X"00",X"06",
		X"10",X"09",X"17",X"02",X"07",X"03",X"1B",X"76",X"C3",X"00",X"00",X"07",X"0E",X"09",X"16",X"01",
		X"08",X"02",X"23",X"77",X"25",X"00",X"00",X"06",X"0A",X"09",X"0A",X"02",X"00",X"02",X"1A",X"77",
		X"61",X"00",X"00",X"06",X"0F",X"09",X"18",X"02",X"09",X"03",X"19",X"77",X"BB",X"00",X"00",X"06",
		X"0C",X"09",X"16",X"01",X"0A",X"03",X"1A",X"78",X"03",X"00",X"00",X"07",X"0D",X"09",X"16",X"01",
		X"09",X"02",X"1A",X"78",X"5E",X"00",X"00",X"07",X"0F",X"09",X"18",X"02",X"09",X"03",X"1A",X"78",
		X"C7",X"00",X"00",X"07",X"0E",X"09",X"17",X"01",X"09",X"03",X"1A",X"79",X"29",X"00",X"00",X"07",
		X"0F",X"09",X"18",X"01",X"09",X"04",X"1A",X"79",X"92",X"00",X"00",X"08",X"0E",X"09",X"17",X"00",
		X"09",X"02",X"23",X"7A",X"02",X"00",X"00",X"05",X"0A",X"09",X"0A",X"02",X"00",X"03",X"26",X"7B",
		X"0A",X"00",X"00",X"07",X"1A",X"09",X"17",X"00",X"FD",X"03",X"23",X"7B",X"C0",X"00",X"00",X"07",
		X"03",X"09",X"03",X"01",X"00",X"03",X"20",X"7B",X"D5",X"00",X"00",X"06",X"05",X"09",X"08",X"01",
		X"03",X"02",X"20",X"7B",X"F3",X"00",X"00",X"06",X"05",X"09",X"08",X"02",X"03",X"03",X"1E",X"7C",
		X"11",X"00",X"00",X"06",X"05",X"09",X"0A",X"01",X"05",X"02",X"1E",X"7C",X"2F",X"00",X"00",X"06",
		X"05",X"09",X"0A",X"02",X"05",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"18",X"95",X"7E",X"1B",X"BC",X"29",X"E0",X"21",X"E8",X"22",X"B4",X"23",X"80",X"24",X"4C",
		X"25",X"18",X"25",X"E4",X"26",X"B0",X"27",X"7C",X"28",X"48",X"29",X"14",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"2A",X"AC",X"0A",X"00",X"00",X"BC",X"9A",X"CD",X"9B",X"0F",X"D0",X"00",
		X"00",X"BC",X"8A",X"CD",X"8B",X"0F",X"D0",X"00",X"00",X"BC",X"7A",X"CD",X"7B",X"0F",X"D0",X"0F",
		X"D0",X"BC",X"8B",X"AB",X"AA",X"CD",X"9B",X"0F",X"D0",X"BC",X"7B",X"AB",X"9A",X"CD",X"8B",X"0F",
		X"D0",X"BC",X"6B",X"AB",X"8A",X"CD",X"7B",X"34",X"70",X"CE",X"18",X"89",X"96",X"49",X"26",X"03",
		X"CE",X"18",X"8F",X"10",X"8E",X"C0",X"01",X"8E",X"C0",X"91",X"8D",X"06",X"8D",X"04",X"8D",X"02",
		X"35",X"F0",X"A6",X"43",X"A7",X"A4",X"A7",X"A9",X"04",X"00",X"A6",X"C0",X"A7",X"84",X"A7",X"89",
		X"04",X"00",X"30",X"88",X"10",X"31",X"A8",X"10",X"39",X"27",X"28",X"29",X"24",X"25",X"26",X"00",
		X"00",X"00",X"24",X"25",X"26",X"34",X"40",X"97",X"BA",X"8E",X"18",X"06",X"3A",X"3A",X"AE",X"84",
		X"9F",X"25",X"BD",X"18",X"57",X"B6",X"18",X"26",X"B7",X"CB",X"40",X"86",X"80",X"B7",X"CB",X"60",
		X"4F",X"5F",X"FD",X"B8",X"14",X"FD",X"91",X"00",X"8E",X"91",X"00",X"ED",X"81",X"ED",X"81",X"ED",
		X"81",X"ED",X"81",X"8C",X"B2",X"EE",X"25",X"F3",X"10",X"8E",X"C0",X"00",X"9E",X"25",X"A6",X"80",
		X"A7",X"A0",X"BD",X"1C",X"12",X"10",X"8C",X"C0",X"60",X"25",X"F3",X"30",X"10",X"C6",X"10",X"A6",
		X"80",X"CE",X"1E",X"1D",X"84",X"7F",X"A6",X"C6",X"6D",X"1F",X"2A",X"02",X"88",X"80",X"A7",X"A0",
		X"34",X"04",X"BD",X"1C",X"12",X"35",X"04",X"5A",X"26",X"E5",X"30",X"88",X"E0",X"10",X"8C",X"C0",
		X"C0",X"25",X"DA",X"BD",X"18",X"57",X"33",X"89",X"00",X"D0",X"10",X"8E",X"D0",X"22",X"E6",X"C4",
		X"C4",X"F0",X"54",X"54",X"54",X"54",X"8E",X"18",X"27",X"3A",X"EC",X"84",X"27",X"0B",X"ED",X"A4",
		X"EC",X"08",X"ED",X"22",X"EC",X"88",X"10",X"ED",X"24",X"E6",X"C0",X"C4",X"0F",X"8E",X"18",X"3F",
		X"3A",X"EC",X"84",X"27",X"0B",X"ED",X"26",X"EC",X"08",X"ED",X"28",X"EC",X"88",X"10",X"ED",X"2A",
		X"31",X"A8",X"20",X"10",X"8C",X"D1",X"20",X"25",X"C5",X"FC",X"18",X"41",X"FD",X"D0",X"5A",X"FC",
		X"18",X"43",X"FD",X"D0",X"5C",X"FC",X"18",X"45",X"FD",X"D0",X"5E",X"CC",X"FF",X"AF",X"FD",X"D0",
		X"22",X"CC",X"BC",X"AC",X"FD",X"D0",X"24",X"CC",X"B1",X"9A",X"FD",X"D0",X"26",X"CC",X"CD",X"7B",
		X"FD",X"D0",X"36",X"CC",X"FF",X"8B",X"FD",X"D0",X"38",X"CC",X"CC",X"AC",X"FD",X"D0",X"3A",X"CC",
		X"CC",X"9C",X"FD",X"D0",X"3C",X"CC",X"CC",X"8C",X"FD",X"D0",X"3E",X"34",X"01",X"1A",X"F0",X"0F",
		X"71",X"86",X"FD",X"97",X"72",X"FC",X"E0",X"9C",X"7D",X"B8",X"14",X"26",X"06",X"BD",X"1B",X"6D",
		X"FC",X"E0",X"86",X"DD",X"6F",X"35",X"01",X"8E",X"91",X"02",X"A6",X"80",X"27",X"FC",X"30",X"1F",
		X"10",X"8E",X"A1",X"02",X"A6",X"A2",X"27",X"FC",X"31",X"A8",X"48",X"10",X"9F",X"62",X"30",X"88",
		X"B8",X"9F",X"60",X"DC",X"62",X"93",X"60",X"DD",X"64",X"CE",X"91",X"02",X"EC",X"81",X"ED",X"C1",
		X"9C",X"62",X"23",X"F8",X"4F",X"5F",X"ED",X"C1",X"11",X"83",X"A3",X"82",X"25",X"F8",X"DC",X"60",
		X"83",X"91",X"02",X"FD",X"91",X"00",X"CC",X"91",X"02",X"DD",X"60",X"DC",X"62",X"B3",X"91",X"00",
		X"DD",X"62",X"8E",X"B7",X"49",X"EC",X"84",X"27",X"16",X"B3",X"91",X"00",X"ED",X"84",X"1F",X"02",
		X"A6",X"A9",X"91",X"02",X"A4",X"02",X"A7",X"02",X"EC",X"03",X"B3",X"91",X"00",X"ED",X"03",X"30",
		X"07",X"8C",X"B7",X"6C",X"23",X"DF",X"10",X"9E",X"64",X"CE",X"FF",X"FA",X"9E",X"60",X"A6",X"80",
		X"85",X"0F",X"27",X"06",X"85",X"10",X"26",X"02",X"33",X"41",X"31",X"3F",X"26",X"F0",X"DF",X"66",
		X"FC",X"B8",X"14",X"26",X"09",X"7C",X"B7",X"48",X"BD",X"E0",X"B3",X"7E",X"1B",X"6B",X"58",X"58",
		X"44",X"56",X"44",X"56",X"B3",X"91",X"00",X"FD",X"B8",X"1B",X"CE",X"91",X"02",X"0F",X"9D",X"8E",
		X"1C",X"02",X"A6",X"C0",X"2F",X"21",X"84",X"0F",X"A6",X"86",X"27",X"1B",X"1F",X"30",X"C3",X"6E",
		X"FD",X"F3",X"91",X"00",X"58",X"49",X"58",X"49",X"54",X"54",X"34",X"02",X"E1",X"E0",X"22",X"07",
		X"0A",X"9D",X"D6",X"9D",X"E7",X"C8",X"BE",X"11",X"93",X"62",X"25",X"D6",X"D6",X"9D",X"50",X"D7",
		X"A4",X"CE",X"91",X"02",X"D6",X"9D",X"8E",X"1C",X"02",X"A6",X"C0",X"2F",X"0F",X"84",X"0F",X"A6",
		X"86",X"27",X"09",X"A6",X"C8",X"BE",X"2B",X"04",X"5A",X"E7",X"C8",X"BE",X"11",X"93",X"62",X"25",
		X"E8",X"50",X"D7",X"9D",X"CE",X"91",X"02",X"10",X"8E",X"B2",X"9A",X"A6",X"C0",X"2C",X"26",X"1F",
		X"30",X"C3",X"6E",X"FD",X"F3",X"91",X"00",X"58",X"49",X"58",X"49",X"54",X"54",X"1E",X"89",X"58",
		X"58",X"44",X"56",X"44",X"56",X"B3",X"91",X"00",X"C3",X"91",X"02",X"1F",X"01",X"A6",X"84",X"E6",
		X"5F",X"40",X"50",X"A7",X"A5",X"11",X"93",X"62",X"25",X"D1",X"CE",X"91",X"02",X"96",X"9D",X"34",
		X"02",X"E6",X"C0",X"2C",X"FC",X"50",X"33",X"C8",X"40",X"8E",X"B8",X"AB",X"3A",X"3A",X"3A",X"3A",
		X"1F",X"12",X"C6",X"01",X"BD",X"1B",X"BC",X"C6",X"02",X"BD",X"1B",X"BC",X"C6",X"04",X"BD",X"1B",
		X"BC",X"C6",X"08",X"BD",X"1B",X"BC",X"33",X"C8",X"C0",X"6A",X"E4",X"26",X"D4",X"35",X"02",X"BE",
		X"B8",X"1B",X"A6",X"89",X"91",X"02",X"84",X"F0",X"A7",X"89",X"91",X"02",X"A6",X"89",X"91",X"42",
		X"84",X"F0",X"A7",X"89",X"91",X"42",X"6F",X"89",X"91",X"82",X"6F",X"89",X"91",X"C2",X"A6",X"89",
		X"92",X"02",X"B7",X"B7",X"46",X"84",X"FD",X"A7",X"89",X"92",X"02",X"31",X"89",X"01",X"00",X"10",
		X"BF",X"B7",X"44",X"A6",X"89",X"91",X"03",X"84",X"F0",X"A7",X"89",X"91",X"03",X"6F",X"89",X"91",
		X"04",X"6F",X"89",X"91",X"05",X"A6",X"89",X"91",X"06",X"B7",X"B7",X"42",X"84",X"FE",X"A7",X"89",
		X"91",X"06",X"31",X"04",X"10",X"BF",X"B7",X"40",X"BD",X"E0",X"93",X"35",X"C0",X"8E",X"1B",X"9C",
		X"10",X"8E",X"D0",X"20",X"EC",X"81",X"27",X"1B",X"ED",X"A4",X"ED",X"A8",X"20",X"ED",X"A8",X"40",
		X"ED",X"A8",X"60",X"ED",X"A9",X"00",X"80",X"ED",X"A9",X"00",X"A0",X"ED",X"A9",X"00",X"C0",X"ED",
		X"A9",X"00",X"E0",X"31",X"22",X"10",X"8C",X"D0",X"40",X"25",X"D9",X"39",X"00",X"00",X"FF",X"DF",
		X"EE",X"C1",X"AE",X"D1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"5F",X"D5",X"0E",X"D1",X"0F",X"90",X"6A",X"DA",X"00",X"00",X"34",X"41",X"1A",X"F0",
		X"1F",X"98",X"A4",X"C4",X"27",X"1B",X"8E",X"1B",X"F0",X"3A",X"3A",X"D7",X"5F",X"EC",X"84",X"33",
		X"CB",X"A6",X"C8",X"BF",X"2B",X"0C",X"8E",X"1B",X"E7",X"D6",X"5F",X"E6",X"85",X"E4",X"C4",X"26",
		X"E5",X"4F",X"40",X"A7",X"A0",X"35",X"C1",X"00",X"07",X"0B",X"00",X"0D",X"00",X"00",X"00",X"0E",
		X"00",X"00",X"FF",X"FF",X"FF",X"C0",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"FF",
		X"FF",X"FF",X"C6",X"0D",X"34",X"76",X"97",X"5F",X"84",X"7F",X"CE",X"1D",X"9D",X"A6",X"C6",X"10",
		X"2B",X"01",X"2B",X"3D",X"CE",X"1E",X"9D",X"33",X"CB",X"31",X"3F",X"1F",X"20",X"58",X"49",X"58",
		X"49",X"58",X"49",X"58",X"49",X"CB",X"0F",X"34",X"06",X"86",X"03",X"3D",X"C3",X"00",X"0C",X"34",
		X"06",X"E6",X"88",X"5F",X"58",X"58",X"E7",X"64",X"54",X"EB",X"88",X"5F",X"4F",X"E3",X"E4",X"ED",
		X"E4",X"E6",X"62",X"86",X"30",X"3D",X"ED",X"62",X"E3",X"E4",X"44",X"56",X"44",X"56",X"44",X"56",
		X"10",X"8E",X"20",X"CC",X"A6",X"AB",X"34",X"02",X"EC",X"61",X"A3",X"63",X"C3",X"02",X"40",X"44",
		X"56",X"44",X"56",X"44",X"56",X"E6",X"AB",X"35",X"02",X"58",X"58",X"44",X"56",X"44",X"56",X"B3",
		X"91",X"00",X"1F",X"01",X"32",X"64",X"10",X"8E",X"20",X"98",X"96",X"5F",X"2A",X"04",X"10",X"8E",
		X"20",X"B2",X"EC",X"A1",X"30",X"8B",X"A6",X"C0",X"27",X"32",X"A6",X"89",X"91",X"02",X"84",X"1F",
		X"10",X"8C",X"20",X"B2",X"23",X"1C",X"34",X"02",X"A6",X"5F",X"84",X"F0",X"AA",X"E4",X"A7",X"E4",
		X"A6",X"5F",X"84",X"05",X"48",X"AA",X"E4",X"A7",X"E4",X"A6",X"5F",X"84",X"0A",X"44",X"AA",X"E0",
		X"20",X"02",X"AA",X"5F",X"84",X"7F",X"AB",X"E4",X"A7",X"89",X"91",X"02",X"A6",X"61",X"34",X"20",
		X"10",X"AE",X"66",X"E6",X"3F",X"C1",X"9D",X"26",X"25",X"81",X"05",X"26",X"21",X"8D",X"71",X"7D",
		X"B8",X"14",X"26",X"62",X"FD",X"B8",X"14",X"31",X"A8",X"EF",X"10",X"BF",X"B8",X"18",X"31",X"A8",
		X"11",X"A6",X"89",X"91",X"02",X"44",X"44",X"84",X"3C",X"B7",X"B8",X"1A",X"20",X"48",X"C1",X"C9",
		X"26",X"12",X"81",X"06",X"26",X"0E",X"8D",X"58",X"25",X"3C",X"34",X"10",X"30",X"01",X"AF",X"A4",
		X"86",X"FE",X"20",X"15",X"C1",X"49",X"26",X"1E",X"81",X"06",X"26",X"1A",X"8D",X"42",X"25",X"26",
		X"34",X"10",X"30",X"88",X"40",X"AF",X"A4",X"86",X"FD",X"A7",X"22",X"EC",X"68",X"C3",X"FF",X"FF",
		X"ED",X"25",X"35",X"10",X"20",X"10",X"C1",X"CC",X"26",X"04",X"81",X"0B",X"27",X"C8",X"C1",X"4C",
		X"26",X"04",X"81",X"0B",X"27",X"D6",X"35",X"20",X"6A",X"61",X"10",X"26",X"FF",X"44",X"35",X"F6",
		X"1F",X"10",X"F3",X"91",X"00",X"34",X"04",X"58",X"49",X"58",X"49",X"35",X"04",X"C4",X"3F",X"39",
		X"34",X"20",X"A6",X"3F",X"2A",X"13",X"1F",X"20",X"C3",X"FF",X"FF",X"C8",X"F0",X"CB",X"C0",X"1F",
		X"02",X"A6",X"3F",X"81",X"00",X"27",X"19",X"20",X"06",X"96",X"BA",X"27",X"13",X"0A",X"BA",X"35",
		X"20",X"10",X"8E",X"B7",X"42",X"31",X"27",X"6D",X"A4",X"26",X"FA",X"AF",X"23",X"1C",X"FE",X"39",
		X"10",X"AE",X"E4",X"6A",X"3F",X"86",X"00",X"A7",X"3E",X"1A",X"01",X"35",X"A0",X"FF",X"00",X"03",
		X"FF",X"FF",X"04",X"06",X"07",X"09",X"0A",X"0B",X"24",X"00",X"01",X"FF",X"04",X"05",X"07",X"00",
		X"01",X"FF",X"0E",X"11",X"12",X"15",X"FF",X"FF",X"FF",X"FF",X"22",X"20",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"16",X"17",X"18",X"16",X"17",X"17",X"18",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1C",X"1E",X"1A",X"1A",X"1A",X"16",X"17",X"18",X"1A",
		X"23",X"1C",X"1F",X"FF",X"FF",X"25",X"25",X"FF",X"26",X"26",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"81",X"82",
		X"83",X"04",X"05",X"86",X"07",X"88",X"89",X"8A",X"0B",X"8C",X"8D",X"8E",X"0F",X"90",X"11",X"92",
		X"93",X"94",X"95",X"96",X"97",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"A0",X"FF",X"FF",
		X"FF",X"29",X"28",X"27",X"26",X"25",X"24",X"2A",X"AB",X"2C",X"AD",X"2E",X"AF",X"B0",X"B1",X"B2",
		X"B3",X"B4",X"35",X"B6",X"B7",X"38",X"39",X"BA",X"BB",X"BC",X"BD",X"BE",X"3F",X"C0",X"41",X"C2",
		X"43",X"C4",X"C5",X"C6",X"C7",X"C8",X"C9",X"CA",X"CB",X"CC",X"CD",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"06",X"02",X"00",X"00",X"04",X"06",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"08",X"00",X"00",
		X"00",X"00",X"04",X"06",X"03",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"09",X"00",X"04",X"06",X"0A",X"00",X"00",X"05",X"06",X"02",X"00",
		X"09",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"0C",X"06",X"02",X"00",X"00",X"04",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"04",X"06",
		X"02",X"00",X"00",X"01",X"00",X"01",X"00",X"09",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"00",
		X"04",X"06",X"03",X"00",X"00",X"00",X"09",X"00",X"04",X"06",X"0A",X"00",X"00",X"05",X"06",X"02",
		X"00",X"09",X"00",X"00",X"00",X"0C",X"06",X"02",X"00",X"00",X"01",X"00",X"01",X"00",X"09",X"00",
		X"09",X"00",X"0C",X"06",X"0A",X"00",X"00",X"05",X"06",X"03",X"00",X"09",X"00",X"09",X"00",X"08",
		X"00",X"08",X"00",X"00",X"24",X"16",X"03",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"08",X"00",
		X"00",X"04",X"06",X"03",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"28",X"00",X"01",X"00",X"19",
		X"00",X"00",X"00",X"2C",X"26",X"22",X"00",X"00",X"00",X"00",X"21",X"00",X"29",X"00",X"00",X"00",
		X"2C",X"16",X"02",X"00",X"00",X"00",X"00",X"00",X"24",X"16",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"19",X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"28",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"24",X"16",X"02",X"00",X"00",X"00",X"00",X"01",X"00",X"09",X"00",X"00",
		X"00",X"0C",X"06",X"02",X"00",X"00",X"00",X"00",X"01",X"00",X"09",X"00",X"04",X"06",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"03",X"00",X"00",X"00",X"09",
		X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"06",X"02",X"00",X"09",X"00",X"08",X"01",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"08",X"00",X"00",X"00",X"00",
		X"04",X"06",X"06",X"06",X"02",X"00",X"00",X"00",X"00",X"01",X"00",X"09",X"00",X"00",X"00",X"0D",
		X"06",X"02",X"00",X"09",X"00",X"08",X"01",X"00",X"09",X"00",X"04",X"06",X"0E",X"06",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"07",X"06",X"02",X"00",X"09",X"00",X"08",
		X"01",X"00",X"09",X"00",X"04",X"06",X"0B",X"00",X"00",X"00",X"09",X"00",X"08",X"01",X"00",X"09",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"02",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"01",X"00",X"09",X"00",X"04",X"06",X"0F",X"06",X"02",X"00",X"09",X"00",
		X"08",X"00",X"05",X"06",X"03",X"00",X"09",X"00",X"09",X"00",X"0C",X"06",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"BF",X"00",X"40",X"00",X"40",
		X"FF",X"3F",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"FF",X"3F",X"00",X"40",X"00",X"40",
		X"FF",X"BF",X"00",X"7E",X"FF",X"BF",X"00",X"01",X"00",X"01",X"FF",X"BD",X"00",X"01",X"00",X"01",
		X"00",X"01",X"00",X"01",X"FF",X"BD",X"00",X"01",X"00",X"01",X"FF",X"BF",X"00",X"00",X"00",X"01",
		X"01",X"01",X"02",X"02",X"02",X"03",X"03",X"03",X"04",X"04",X"04",X"05",X"05",X"05",X"06",X"06",
		X"06",X"07",X"07",X"07",X"08",X"08",X"08",X"09",X"09",X"09",X"0A",X"0A",X"0A",X"0B",X"0B",X"0B",
		X"0C",X"0C",X"0C",X"0D",X"0D",X"0D",X"0E",X"0E",X"0E",X"0F",X"0F",X"0F",X"10",X"10",X"10",X"11",
		X"11",X"11",X"12",X"12",X"12",X"13",X"13",X"13",X"14",X"14",X"14",X"15",X"15",X"15",X"16",X"16",
		X"16",X"17",X"17",X"17",X"18",X"18",X"18",X"19",X"19",X"19",X"1A",X"1A",X"1A",X"1B",X"1B",X"1B",
		X"1C",X"1C",X"1C",X"1D",X"1D",X"1D",X"1E",X"1E",X"1E",X"1F",X"1F",X"1F",X"20",X"20",X"20",X"21",
		X"21",X"21",X"22",X"22",X"22",X"23",X"23",X"23",X"24",X"24",X"24",X"25",X"25",X"25",X"26",X"26",
		X"26",X"27",X"27",X"27",X"28",X"28",X"28",X"29",X"29",X"29",X"2A",X"2A",X"2A",X"2B",X"2B",X"2B",
		X"2C",X"2C",X"2C",X"2D",X"2D",X"2D",X"2E",X"2E",X"2E",X"2F",X"2F",X"2F",X"30",X"30",X"30",X"31",
		X"31",X"31",X"32",X"32",X"32",X"33",X"33",X"33",X"34",X"34",X"34",X"35",X"35",X"35",X"36",X"36",
		X"36",X"37",X"37",X"37",X"38",X"38",X"38",X"39",X"39",X"39",X"3A",X"3A",X"3A",X"3B",X"3B",X"3B",
		X"3C",X"3C",X"3C",X"3D",X"3D",X"3D",X"3E",X"3E",X"3E",X"3F",X"3F",X"3F",X"40",X"40",X"40",X"41",
		X"41",X"41",X"42",X"42",X"42",X"43",X"43",X"43",X"44",X"44",X"44",X"45",X"45",X"45",X"46",X"46",
		X"46",X"47",X"47",X"47",X"48",X"48",X"48",X"49",X"49",X"49",X"4A",X"4A",X"4A",X"4B",X"4B",X"4B",
		X"4C",X"4C",X"4C",X"4D",X"4D",X"4D",X"4E",X"4E",X"4E",X"4F",X"4F",X"4F",X"50",X"50",X"50",X"51",
		X"51",X"51",X"52",X"52",X"52",X"53",X"53",X"53",X"54",X"54",X"54",X"55",X"55",X"55",X"56",X"56",
		X"56",X"57",X"57",X"57",X"58",X"58",X"58",X"59",X"59",X"59",X"5A",X"5A",X"5A",X"5B",X"5B",X"5B",
		X"5C",X"5C",X"5C",X"5D",X"26",X"2C",X"2C",X"26",X"00",X"24",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"00",X"00",X"00",X"46",X"C0",X"C7",
		X"01",X"04",X"01",X"18",X"C7",X"00",X"00",X"00",X"00",X"26",X"00",X"00",X"46",X"3C",X"3D",X"15",
		X"07",X"01",X"93",X"42",X"C2",X"C7",X"00",X"00",X"00",X"00",X"00",X"46",X"3C",X"3D",X"12",X"89",
		X"89",X"93",X"44",X"B4",X"3C",X"C5",X"C7",X"00",X"00",X"00",X"46",X"44",X"3D",X"12",X"08",X"08",
		X"16",X"44",X"34",X"C4",X"3D",X"33",X"41",X"00",X"00",X"1D",X"1E",X"36",X"12",X"89",X"06",X"93",
		X"42",X"36",X"C2",X"37",X"C2",X"3C",X"41",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"08",
		X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"08",X"08",
		X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"22",X"22",X"24",X"24",X"24",X"24",
		X"26",X"2C",X"2C",X"26",X"00",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"83",X"83",X"00",X"83",
		X"00",X"00",X"00",X"00",X"00",X"25",X"00",X"46",X"C0",X"B6",X"C0",X"C0",X"95",X"0A",X"86",X"0B",
		X"82",X"00",X"00",X"00",X"00",X"26",X"46",X"3C",X"3E",X"43",X"35",X"3A",X"41",X"05",X"0A",X"0F",
		X"93",X"C0",X"C7",X"00",X"00",X"00",X"3F",X"3E",X"35",X"3E",X"2E",X"45",X"15",X"08",X"08",X"93",
		X"44",X"BE",X"41",X"00",X"00",X"00",X"38",X"43",X"3E",X"3E",X"3D",X"12",X"08",X"08",X"16",X"3C",
		X"BE",X"BA",X"41",X"00",X"00",X"1D",X"1E",X"36",X"2F",X"3D",X"15",X"8A",X"08",X"16",X"44",X"31",
		X"BC",X"BE",X"41",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"08",
		X"08",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"08",
		X"08",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"08",
		X"08",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"02",X"22",X"22",X"22",X"24",X"24",X"24",X"22",X"2C",X"2C",X"22",
		X"00",X"24",X"00",X"00",X"4A",X"49",X"C7",X"00",X"00",X"00",X"00",X"83",X"46",X"C7",X"00",X"00",
		X"00",X"25",X"00",X"46",X"B6",X"42",X"15",X"82",X"4D",X"4C",X"86",X"16",X"3C",X"C5",X"C7",X"00",
		X"00",X"26",X"46",X"44",X"BA",X"2A",X"8A",X"90",X"82",X"01",X"16",X"3C",X"43",X"35",X"41",X"00",
		X"00",X"46",X"B0",X"3E",X"45",X"15",X"89",X"11",X"89",X"16",X"B0",X"BA",X"35",X"43",X"39",X"00",
		X"00",X"C6",X"C4",X"B2",X"12",X"08",X"09",X"0F",X"16",X"44",X"35",X"3B",X"BA",X"3E",X"41",X"00",
		X"00",X"1D",X"1E",X"47",X"81",X"10",X"0B",X"93",X"44",X"35",X"43",X"35",X"43",X"BA",X"39",X"00",
		X"10",X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"22",X"24",X"24",X"24",X"24",X"24",X"1F",X"2E",X"2E",X"1F",X"00",X"24",X"00",X"00",
		X"00",X"00",X"46",X"C7",X"00",X"46",X"C7",X"46",X"C7",X"00",X"00",X"00",X"00",X"25",X"00",X"00",
		X"4A",X"49",X"42",X"12",X"0C",X"96",X"C2",X"3C",X"32",X"C7",X"00",X"00",X"00",X"26",X"00",X"46",
		X"B6",X"42",X"15",X"08",X"08",X"09",X"96",X"C4",X"3E",X"32",X"C7",X"00",X"00",X"00",X"46",X"B3",
		X"45",X"12",X"89",X"88",X"88",X"10",X"89",X"96",X"C4",X"3E",X"41",X"00",X"00",X"00",X"38",X"45",
		X"15",X"08",X"08",X"89",X"09",X"88",X"09",X"0F",X"96",X"C4",X"39",X"00",X"00",X"1D",X"1E",X"47",
		X"81",X"88",X"08",X"08",X"89",X"88",X"10",X"02",X"05",X"96",X"47",X"00",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",
		X"10",X"10",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",
		X"10",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"22",X"22",X"22",X"22",
		X"24",X"24",X"24",X"24",X"1F",X"29",X"29",X"1F",X"00",X"24",X"00",X"00",X"4A",X"49",X"C7",X"46",
		X"B6",X"B6",X"C7",X"01",X"0E",X"00",X"00",X"00",X"00",X"25",X"00",X"00",X"46",X"3C",X"BD",X"AF",
		X"BA",X"45",X"12",X"08",X"08",X"0E",X"00",X"00",X"00",X"26",X"00",X"46",X"3C",X"3E",X"2D",X"3E",
		X"3D",X"15",X"89",X"89",X"89",X"89",X"04",X"00",X"00",X"00",X"46",X"3C",X"2C",X"2C",X"2D",X"3A",
		X"2A",X"11",X"11",X"11",X"11",X"07",X"00",X"00",X"00",X"00",X"3F",X"3E",X"2D",X"3E",X"3A",X"2D",
		X"C5",X"95",X"09",X"09",X"09",X"09",X"04",X"00",X"00",X"1D",X"1E",X"30",X"43",X"3A",X"BE",X"2D",
		X"3E",X"C5",X"92",X"88",X"88",X"8E",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"1E",X"2E",X"2E",X"1E",X"00",X"24",X"00",X"00",X"00",X"83",X"46",X"C7",X"46",X"B6",X"C7",X"46",
		X"B6",X"C7",X"00",X"00",X"00",X"25",X"00",X"00",X"01",X"90",X"96",X"C2",X"42",X"C4",X"C5",X"42",
		X"C4",X"C5",X"C7",X"00",X"00",X"26",X"46",X"C0",X"95",X"88",X"88",X"96",X"C2",X"42",X"C4",X"C5",
		X"42",X"C4",X"39",X"00",X"00",X"00",X"3F",X"3E",X"41",X"05",X"08",X"90",X"96",X"C2",X"42",X"C4",
		X"C5",X"42",X"47",X"00",X"00",X"00",X"38",X"45",X"15",X"08",X"08",X"0A",X"88",X"96",X"C2",X"42",
		X"C4",X"C5",X"C7",X"00",X"00",X"1D",X"1E",X"47",X"81",X"8A",X"02",X"81",X"10",X"16",X"42",X"C2",
		X"42",X"C4",X"39",X"00",X"10",X"10",X"10",X"10",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"22",X"22",X"24",X"24",X"24",X"24",X"24",X"21",X"2D",X"2D",X"21",
		X"00",X"24",X"00",X"00",X"4A",X"49",X"B6",X"C7",X"46",X"B6",X"B6",X"C7",X"83",X"00",X"00",X"00",
		X"00",X"25",X"00",X"00",X"00",X"38",X"BB",X"32",X"3C",X"3E",X"3D",X"15",X"90",X"82",X"00",X"00",
		X"00",X"26",X"00",X"00",X"46",X"3C",X"3E",X"3E",X"BB",X"45",X"15",X"89",X"06",X"0A",X"82",X"00",
		X"00",X"00",X"00",X"46",X"3C",X"3E",X"3E",X"BB",X"45",X"12",X"06",X"09",X"86",X"8A",X"02",X"00",
		X"00",X"00",X"46",X"3C",X"3E",X"3E",X"BB",X"45",X"15",X"90",X"82",X"81",X"10",X"06",X"04",X"00",
		X"00",X"1D",X"1E",X"33",X"BB",X"BB",X"45",X"15",X"89",X"06",X"0A",X"82",X"81",X"04",X"00",X"00",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"25",X"2B",X"2B",X"25",X"00",X"24",X"00",X"00",
		X"4A",X"49",X"B6",X"C7",X"83",X"83",X"00",X"46",X"C7",X"00",X"00",X"00",X"00",X"25",X"00",X"46",
		X"C0",X"B3",X"45",X"15",X"06",X"07",X"46",X"B0",X"C5",X"C7",X"00",X"00",X"00",X"26",X"46",X"B0",
		X"35",X"45",X"15",X"02",X"01",X"16",X"44",X"AD",X"3D",X"15",X"04",X"00",X"00",X"46",X"B0",X"35",
		X"45",X"15",X"06",X"86",X"16",X"44",X"AD",X"3D",X"15",X"07",X"00",X"00",X"00",X"C6",X"33",X"45",
		X"15",X"02",X"01",X"16",X"44",X"AD",X"3D",X"15",X"8A",X"89",X"04",X"00",X"00",X"1D",X"1E",X"47",
		X"81",X"86",X"16",X"44",X"AD",X"3D",X"15",X"0B",X"0B",X"07",X"00",X"00",X"18",X"18",X"18",X"18",
		X"18",X"18",X"18",X"10",X"10",X"10",X"10",X"08",X"08",X"00",X"00",X"00",X"18",X"18",X"18",X"18",
		X"18",X"18",X"18",X"10",X"10",X"10",X"10",X"08",X"08",X"00",X"00",X"00",X"18",X"18",X"18",X"18",
		X"18",X"18",X"10",X"10",X"10",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"18",X"18",X"18",X"18",
		X"18",X"10",X"10",X"10",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"18",X"18",X"18",X"18",
		X"10",X"10",X"10",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"18",X"18",
		X"10",X"10",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"22",X"22",
		X"22",X"42",X"42",X"42",X"1E",X"2A",X"2A",X"1E",X"00",X"24",X"00",X"46",X"B6",X"C7",X"83",X"46",
		X"B6",X"B6",X"B6",X"B6",X"C7",X"00",X"00",X"00",X"00",X"25",X"46",X"B3",X"45",X"C2",X"95",X"13",
		X"C4",X"BA",X"2D",X"BB",X"C5",X"C7",X"00",X"00",X"00",X"26",X"38",X"BB",X"B1",X"AF",X"BD",X"92",
		X"96",X"BC",X"43",X"AD",X"2D",X"BD",X"C7",X"00",X"00",X"00",X"38",X"3B",X"B2",X"30",X"3D",X"12",
		X"93",X"3C",X"BB",X"43",X"2C",X"45",X"47",X"00",X"00",X"00",X"38",X"3E",X"C5",X"42",X"15",X"90",
		X"96",X"C4",X"AD",X"3B",X"43",X"39",X"00",X"00",X"00",X"1D",X"1E",X"36",X"36",X"12",X"89",X"0B",
		X"0A",X"96",X"BC",X"3A",X"AD",X"C5",X"C7",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"08",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"08",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"22",X"22",X"24",X"24",X"24",X"24",
		X"23",X"2B",X"2B",X"23",X"00",X"24",X"00",X"00",X"46",X"B6",X"C7",X"00",X"00",X"83",X"00",X"83",
		X"00",X"00",X"00",X"00",X"00",X"25",X"00",X"46",X"B3",X"43",X"B1",X"C0",X"97",X"06",X"86",X"8A",
		X"0C",X"82",X"00",X"00",X"00",X"26",X"46",X"B3",X"43",X"3E",X"3E",X"2C",X"BD",X"97",X"06",X"89",
		X"90",X"0B",X"04",X"00",X"00",X"00",X"38",X"43",X"3E",X"43",X"AD",X"43",X"2D",X"C5",X"97",X"06",
		X"8A",X"8A",X"04",X"00",X"00",X"00",X"38",X"3A",X"3D",X"2B",X"BC",X"2E",X"3E",X"B2",X"C2",X"97",
		X"8D",X"89",X"04",X"00",X"00",X"1D",X"1E",X"36",X"12",X"0B",X"96",X"C4",X"31",X"C2",X"B0",X"BD",
		X"97",X"89",X"04",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",
		X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"10",X"10",X"08",X"08",X"08",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"22",X"22",X"22",X"22",X"42",X"42",X"42",X"42",X"1E",X"2A",X"2A",X"1E",
		X"00",X"24",X"00",X"00",X"00",X"00",X"46",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"C7",X"00",X"00",
		X"00",X"25",X"00",X"00",X"00",X"46",X"44",X"43",X"43",X"43",X"43",X"43",X"43",X"C5",X"C7",X"00",
		X"00",X"26",X"00",X"00",X"46",X"44",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"39",X"00",
		X"00",X"00",X"00",X"46",X"44",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"39",X"00",
		X"00",X"00",X"46",X"44",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"39",X"00",
		X"00",X"46",X"44",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"39",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"15",X"1D",X"1D",X"15",X"00",X"24",X"00",X"00",
		X"4A",X"49",X"B6",X"C7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"00",X"46",
		X"B6",X"44",X"45",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"26",X"46",X"B3",
		X"43",X"45",X"15",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"43",
		X"45",X"15",X"0B",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"45",
		X"15",X"06",X"0B",X"0B",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1D",X"1E",X"47",
		X"03",X"00",X"05",X"0B",X"0B",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",
		X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"30",X"D4",X"30",X"EB",X"31",X"02",X"31",X"19",X"31",X"30",X"31",X"47",X"31",X"5E",X"31",X"75",
		X"31",X"8C",X"31",X"A3",X"31",X"BA",X"31",X"BF",X"31",X"D6",X"31",X"ED",X"32",X"04",X"32",X"1B",
		X"32",X"32",X"32",X"49",X"32",X"60",X"32",X"77",X"32",X"87",X"32",X"9E",X"32",X"B5",X"32",X"CC",
		X"32",X"EA",X"33",X"01",X"33",X"18",X"33",X"2F",X"33",X"46",X"33",X"5D",X"33",X"74",X"33",X"8B",
		X"33",X"A2",X"33",X"B9",X"33",X"D7",X"33",X"EE",X"34",X"05",X"34",X"1C",X"34",X"33",X"34",X"3F",
		X"34",X"49",X"34",X"60",X"34",X"70",X"34",X"80",X"34",X"90",X"34",X"96",X"34",X"A8",X"34",X"B1",
		X"34",X"CF",X"34",X"E6",X"34",X"EE",X"34",X"F5",X"35",X"0F",X"35",X"26",X"35",X"32",X"35",X"3E",
		X"35",X"4A",X"35",X"56",X"35",X"62",X"35",X"6E",X"35",X"7A",X"35",X"86",X"35",X"92",X"35",X"9E",
		X"35",X"AA",X"35",X"B6",X"35",X"C2",X"35",X"CE",X"35",X"DA",X"35",X"E6",X"35",X"F2",X"35",X"FE",
		X"36",X"0A",X"36",X"16",X"36",X"22",X"36",X"2E",X"36",X"3A",X"36",X"4B",X"35",X"26",X"36",X"57",
		X"36",X"63",X"36",X"6F",X"35",X"62",X"36",X"7B",X"36",X"87",X"36",X"93",X"36",X"9F",X"36",X"B0",
		X"36",X"BC",X"36",X"C8",X"36",X"D4",X"36",X"E0",X"36",X"EA",X"36",X"F2",X"36",X"FE",X"37",X"05",
		X"37",X"11",X"37",X"1D",X"37",X"21",X"37",X"28",X"37",X"2F",X"37",X"40",X"37",X"60",X"37",X"28",
		X"37",X"28",X"37",X"28",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"10",X"01",X"10",X"10",
		X"10",X"10",X"11",X"00",X"10",X"10",X"00",X"10",X"01",X"11",X"00",X"03",X"07",X"00",X"10",X"00",
		X"01",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"11",
		X"11",X"10",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"00",X"00",X"10",X"00",X"11",X"00",
		X"01",X"00",X"00",X"10",X"00",X"10",X"11",X"11",X"10",X"03",X"07",X"01",X"11",X"00",X"10",X"00",
		X"10",X"00",X"00",X"10",X"00",X"11",X"00",X"00",X"00",X"10",X"10",X"00",X"10",X"01",X"11",X"00",
		X"03",X"07",X"00",X"01",X"10",X"00",X"10",X"10",X"01",X"00",X"10",X"10",X"00",X"10",X"11",X"11",
		X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"03",X"07",X"11",X"11",X"10",X"10",X"00",X"00",X"11",
		X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"10",X"00",X"10",X"01",X"11",X"00",X"03",X"07",
		X"01",X"11",X"00",X"10",X"00",X"00",X"10",X"11",X"00",X"11",X"00",X"10",X"10",X"00",X"10",X"10",
		X"00",X"10",X"01",X"11",X"00",X"03",X"07",X"11",X"11",X"10",X"10",X"00",X"10",X"00",X"01",X"00",
		X"00",X"10",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"03",X"07",X"01",X"11",
		X"00",X"10",X"00",X"10",X"10",X"00",X"10",X"01",X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"10",
		X"01",X"11",X"00",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"10",X"10",X"01",
		X"10",X"01",X"10",X"10",X"00",X"00",X"10",X"01",X"11",X"00",X"03",X"01",X"00",X"00",X"00",X"03",
		X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"10",X"11",X"11",X"10",X"10",X"00",X"10",
		X"10",X"00",X"10",X"10",X"00",X"10",X"03",X"07",X"11",X"11",X"00",X"10",X"00",X"10",X"10",X"00",
		X"10",X"10",X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"10",X"11",X"11",X"00",X"03",X"07",X"01",
		X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",
		X"10",X"01",X"11",X"00",X"03",X"07",X"11",X"10",X"00",X"10",X"01",X"00",X"10",X"00",X"10",X"10",
		X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"11",X"11",X"00",X"03",X"07",X"01",X"11",X"00",
		X"10",X"00",X"10",X"10",X"00",X"00",X"11",X"11",X"00",X"10",X"00",X"00",X"10",X"00",X"10",X"01",
		X"11",X"00",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"00",X"11",X"11",X"00",
		X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"03",X"07",X"01",X"11",X"00",X"10",X"00",
		X"10",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"01",X"10",X"10",X"00",X"10",X"01",X"11",X"00",
		X"03",X"07",X"01",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"11",X"11",X"10",X"10",X"00",
		X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"02",X"07",X"11",X"10",X"01",X"00",X"01",X"00",X"01",
		X"00",X"01",X"00",X"01",X"00",X"11",X"10",X"03",X"07",X"00",X"01",X"10",X"00",X"00",X"10",X"00",
		X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"10",X"00",X"10",X"01",X"11",X"00",X"03",X"07",
		X"10",X"00",X"10",X"10",X"01",X"00",X"10",X"10",X"00",X"11",X"00",X"00",X"10",X"10",X"00",X"10",
		X"01",X"00",X"10",X"00",X"10",X"03",X"07",X"01",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",
		X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"10",X"11",X"11",X"10",X"04",X"07",X"01",X"10",
		X"11",X"00",X"10",X"01",X"00",X"10",X"10",X"01",X"00",X"10",X"10",X"01",X"00",X"10",X"10",X"01",
		X"00",X"10",X"10",X"00",X"00",X"10",X"01",X"00",X"01",X"00",X"03",X"07",X"10",X"00",X"10",X"11",
		X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"01",X"10",X"10",X"00",
		X"10",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"10",
		X"00",X"10",X"10",X"00",X"10",X"01",X"11",X"00",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",
		X"10",X"00",X"10",X"11",X"11",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"03",
		X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"10",X"10",X"10",
		X"10",X"01",X"00",X"01",X"10",X"10",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"10",X"00",
		X"10",X"11",X"11",X"00",X"10",X"10",X"00",X"10",X"01",X"00",X"10",X"00",X"10",X"03",X"07",X"01",
		X"11",X"00",X"10",X"00",X"10",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"10",X"00",
		X"10",X"01",X"11",X"00",X"03",X"07",X"01",X"11",X"00",X"10",X"10",X"10",X"00",X"10",X"00",X"00",
		X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"01",X"11",X"00",X"03",X"07",X"01",X"00",X"10",
		X"10",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"01",
		X"11",X"00",X"03",X"07",X"01",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",
		X"01",X"01",X"00",X"01",X"01",X"00",X"00",X"10",X"00",X"04",X"07",X"01",X"00",X"01",X"00",X"10",
		X"00",X"00",X"10",X"10",X"00",X"00",X"10",X"10",X"01",X"00",X"10",X"10",X"01",X"00",X"10",X"10",
		X"01",X"00",X"10",X"01",X"10",X"11",X"00",X"03",X"07",X"10",X"00",X"10",X"10",X"00",X"10",X"01",
		X"01",X"00",X"00",X"10",X"00",X"01",X"01",X"00",X"10",X"00",X"10",X"10",X"00",X"10",X"03",X"07",
		X"01",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"01",X"01",X"00",X"00",X"10",X"00",X"00",
		X"10",X"00",X"00",X"10",X"00",X"03",X"07",X"01",X"11",X"10",X"00",X"00",X"10",X"00",X"01",X"00",
		X"00",X"10",X"00",X"01",X"00",X"00",X"10",X"00",X"00",X"11",X"11",X"10",X"03",X"07",X"00",X"0A",
		X"00",X"00",X"A0",X"00",X"0A",X"00",X"00",X"AA",X"AA",X"A0",X"0A",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"0A",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"AA",X"B0",X"00",X"00",X"AA",X"B0",X"02",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"B0",X"03",X"07",X"0A",X"AB",X"00",X"AA",X"BA",
		X"B0",X"AB",X"0A",X"B0",X"00",X"AB",X"00",X"0A",X"B0",X"00",X"00",X"00",X"00",X"0A",X"B0",X"00",
		X"02",X"07",X"0A",X"B0",X"AA",X"B0",X"0A",X"B0",X"0A",X"B0",X"0A",X"B0",X"00",X"00",X"0A",X"B0",
		X"02",X"07",X"0A",X"B0",X"AA",X"B0",X"AB",X"00",X"AB",X"00",X"AB",X"00",X"AA",X"B0",X"0A",X"B0",
		X"02",X"07",X"AB",X"00",X"AA",X"B0",X"0A",X"B0",X"0A",X"B0",X"0A",X"B0",X"AA",X"B0",X"AB",X"00",
		X"02",X"02",X"AA",X"B0",X"AB",X"00",X"02",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"A0",X"0A",X"A0",X"A0",X"00",X"01",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"03",X"07",X"00",X"00",X"AA",X"00",X"00",X"00",X"AB",X"00",X"00",X"0A",X"B0",X"00",X"00",
		X"AB",X"00",X"00",X"0A",X"B0",X"00",X"00",X"AB",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"03",
		X"07",X"0A",X"00",X"00",X"A0",X"A0",X"00",X"A0",X"A0",X"00",X"0A",X"00",X"00",X"A0",X"A0",X"A0",
		X"A0",X"0A",X"00",X"0A",X"A0",X"A0",X"03",X"02",X"AA",X"0A",X"A0",X"AB",X"0A",X"B0",X"01",X"05",
		X"00",X"00",X"A0",X"00",X"A0",X"03",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"A0",X"03",
		X"07",X"00",X"A0",X"00",X"0A",X"AA",X"00",X"A0",X"A0",X"A0",X"00",X"A0",X"00",X"00",X"A0",X"00",
		X"00",X"A0",X"00",X"00",X"A0",X"00",X"02",X"05",X"AA",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"AA",X"A0",X"02",X"05",X"0A",X"00",X"AA",X"00",X"0A",X"00",X"0A",X"00",X"AA",X"A0",X"02",X"05",
		X"AA",X"A0",X"00",X"A0",X"AA",X"A0",X"A0",X"00",X"AA",X"A0",X"02",X"05",X"AA",X"A0",X"00",X"A0",
		X"AA",X"A0",X"00",X"A0",X"AA",X"A0",X"02",X"05",X"A0",X"A0",X"A0",X"A0",X"AA",X"A0",X"00",X"A0",
		X"00",X"A0",X"02",X"05",X"AA",X"A0",X"A0",X"00",X"AA",X"A0",X"00",X"A0",X"AA",X"A0",X"02",X"05",
		X"AA",X"A0",X"A0",X"00",X"AA",X"A0",X"A0",X"A0",X"AA",X"A0",X"02",X"05",X"AA",X"A0",X"00",X"A0",
		X"0A",X"00",X"0A",X"00",X"0A",X"00",X"02",X"05",X"AA",X"A0",X"A0",X"A0",X"AA",X"A0",X"A0",X"A0",
		X"AA",X"A0",X"02",X"05",X"AA",X"A0",X"A0",X"A0",X"AA",X"A0",X"00",X"A0",X"00",X"A0",X"02",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"AA",X"A0",X"A0",X"A0",
		X"AA",X"A0",X"A0",X"A0",X"A0",X"A0",X"02",X"05",X"AA",X"A0",X"A0",X"A0",X"AA",X"00",X"A0",X"A0",
		X"AA",X"A0",X"02",X"05",X"AA",X"A0",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"AA",X"A0",X"02",X"05",
		X"AA",X"00",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"AA",X"00",X"02",X"05",X"AA",X"A0",X"A0",X"00",
		X"AA",X"00",X"A0",X"00",X"AA",X"A0",X"02",X"05",X"AA",X"A0",X"A0",X"00",X"AA",X"00",X"A0",X"00",
		X"A0",X"00",X"02",X"05",X"AA",X"A0",X"A0",X"00",X"A0",X"A0",X"A0",X"A0",X"AA",X"A0",X"02",X"05",
		X"A0",X"A0",X"A0",X"A0",X"AA",X"A0",X"A0",X"A0",X"A0",X"A0",X"02",X"05",X"AA",X"A0",X"0A",X"00",
		X"0A",X"00",X"0A",X"00",X"AA",X"A0",X"02",X"05",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"A0",X"A0",
		X"AA",X"A0",X"02",X"05",X"A0",X"A0",X"A0",X"A0",X"AA",X"00",X"A0",X"A0",X"A0",X"A0",X"02",X"05",
		X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"AA",X"A0",X"03",X"05",X"AA",X"AA",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"00",X"A0",X"A0",X"00",X"A0",X"02",X"05",X"AA",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"02",X"05",X"AA",X"A0",X"A0",X"A0",X"AA",X"A0",X"A0",
		X"00",X"A0",X"00",X"02",X"05",X"AA",X"A0",X"A0",X"A0",X"A0",X"A0",X"0A",X"00",X"00",X"A0",X"02",
		X"05",X"AA",X"A0",X"A0",X"A0",X"AA",X"00",X"A0",X"A0",X"A0",X"A0",X"02",X"05",X"AA",X"A0",X"0A",
		X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"02",X"05",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"AA",X"A0",X"02",X"05",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"0A",X"00",X"0A",X"00",X"03",
		X"05",X"A0",X"00",X"A0",X"A0",X"00",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"AA",X"AA",X"A0",
		X"02",X"05",X"A0",X"A0",X"A0",X"A0",X"0A",X"00",X"A0",X"A0",X"A0",X"A0",X"02",X"05",X"A0",X"A0",
		X"A0",X"A0",X"AA",X"A0",X"0A",X"00",X"0A",X"00",X"02",X"05",X"AA",X"A0",X"00",X"A0",X"0A",X"00",
		X"A0",X"00",X"AA",X"A0",X"02",X"05",X"00",X"A0",X"0A",X"00",X"AA",X"A0",X"0A",X"00",X"00",X"A0",
		X"02",X"04",X"00",X"00",X"AA",X"A0",X"00",X"00",X"AA",X"A0",X"02",X"03",X"00",X"00",X"00",X"00",
		X"AA",X"A0",X"02",X"05",X"AA",X"A0",X"00",X"A0",X"0A",X"A0",X"00",X"00",X"0A",X"00",X"01",X"05",
		X"A0",X"A0",X"A0",X"00",X"A0",X"02",X"05",X"00",X"A0",X"0A",X"00",X"A0",X"00",X"0A",X"00",X"00",
		X"A0",X"02",X"05",X"A0",X"00",X"0A",X"00",X"00",X"A0",X"0A",X"00",X"A0",X"00",X"01",X"02",X"A0",
		X"A0",X"01",X"05",X"00",X"00",X"00",X"A0",X"A0",X"01",X"05",X"00",X"00",X"00",X"00",X"A0",X"03",
		X"05",X"00",X"00",X"A0",X"00",X"0A",X"00",X"00",X"A0",X"00",X"0A",X"00",X"00",X"A0",X"00",X"00",
		X"06",X"05",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",
		X"03",X"05",X"00",X"A0",X"00",X"00",X"0A",X"00",X"AA",X"AA",X"A0",X"00",X"0A",X"00",X"00",X"A0",
		X"00",X"20",X"49",X"4E",X"46",X"45",X"52",X"4E",X"4F",X"20",X"2D",X"20",X"28",X"43",X"29",X"31",
		X"39",X"38",X"34",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"48",X"7E",X"21",X"0F",X"21",X"0F",X"21",X"0F",X"31",X"0F",X"31",X"0F",X"31",X"0F",X"31",
		X"0F",X"31",X"0F",X"41",X"00",X"31",X"0F",X"31",X"0F",X"31",X"0F",X"41",X"0F",X"41",X"0F",X"41",
		X"0F",X"41",X"0F",X"41",X"0F",X"51",X"0F",X"51",X"0F",X"51",X"0F",X"51",X"0F",X"51",X"0F",X"51",
		X"0F",X"51",X"0F",X"51",X"0F",X"51",X"0F",X"61",X"0F",X"61",X"0F",X"61",X"0F",X"61",X"0F",X"61",
		X"0F",X"61",X"20",X"12",X"0F",X"61",X"00",X"51",X"0F",X"51",X"20",X"12",X"0F",X"61",X"0F",X"61",
		X"0F",X"61",X"0F",X"61",X"20",X"12",X"0F",X"61",X"20",X"12",X"0F",X"61",X"0F",X"71",X"0F",X"71",
		X"20",X"12",X"0F",X"71",X"20",X"12",X"0F",X"71",X"20",X"12",X"0F",X"71",X"20",X"12",X"0F",X"71",
		X"20",X"12",X"0F",X"71",X"20",X"22",X"0F",X"81",X"10",X"22",X"0F",X"81",X"20",X"12",X"0F",X"81",
		X"20",X"12",X"0F",X"81",X"20",X"22",X"0F",X"81",X"20",X"22",X"0F",X"91",X"10",X"22",X"0F",X"91",
		X"20",X"12",X"0F",X"91",X"20",X"12",X"0F",X"91",X"20",X"22",X"0F",X"A1",X"10",X"22",X"0F",X"A1",
		X"20",X"12",X"0F",X"A1",X"20",X"12",X"0F",X"A1",X"20",X"12",X"0F",X"A1",X"20",X"22",X"0F",X"B1",
		X"10",X"22",X"0F",X"B1",X"20",X"12",X"0F",X"B1",X"20",X"12",X"0F",X"B1",X"20",X"12",X"0F",X"B1",
		X"20",X"22",X"0F",X"C1",X"10",X"22",X"0F",X"C1",X"20",X"12",X"0F",X"C1",X"20",X"12",X"0F",X"C1",
		X"20",X"12",X"0F",X"C1",X"20",X"22",X"0F",X"C1",X"20",X"22",X"0F",X"C1",X"20",X"22",X"0F",X"D1",
		X"10",X"22",X"0F",X"D1",X"20",X"12",X"0F",X"D1",X"20",X"22",X"0F",X"D1",X"20",X"22",X"0F",X"D1",
		X"20",X"22",X"0F",X"D1",X"20",X"22",X"0F",X"D1",X"20",X"22",X"0F",X"D1",X"20",X"32",X"0F",X"E1",
		X"10",X"32",X"0F",X"E1",X"20",X"22",X"0F",X"E1",X"20",X"22",X"0F",X"E1",X"20",X"22",X"0F",X"E1",
		X"20",X"32",X"00",X"F0",X"42",X"00",X"E2",X"10",X"42",X"00",X"E2",X"10",X"42",X"00",X"E2",X"10",
		X"42",X"00",X"E2",X"10",X"42",X"00",X"E2",X"10",X"42",X"00",X"E2",X"10",X"42",X"00",X"E2",X"10",
		X"42",X"00",X"E2",X"10",X"42",X"00",X"E2",X"10",X"42",X"00",X"E2",X"10",X"42",X"00",X"E2",X"10",
		X"42",X"00",X"E2",X"10",X"42",X"00",X"E2",X"10",X"42",X"00",X"E2",X"10",X"42",X"00",X"E2",X"10",
		X"32",X"00",X"E2",X"10",X"32",X"00",X"E2",X"10",X"22",X"00",X"E2",X"10",X"22",X"00",X"E2",X"10",
		X"12",X"00",X"E2",X"10",X"12",X"FF",X"41",X"30",X"31",X"0F",X"41",X"40",X"21",X"0F",X"41",X"40",
		X"21",X"0F",X"51",X"10",X"12",X"20",X"21",X"0F",X"51",X"40",X"21",X"00",X"41",X"20",X"12",X"10",
		X"31",X"0F",X"51",X"10",X"12",X"20",X"21",X"0F",X"51",X"20",X"12",X"10",X"31",X"0F",X"51",X"20",
		X"12",X"20",X"21",X"0F",X"61",X"10",X"12",X"20",X"31",X"00",X"51",X"20",X"12",X"10",X"31",X"0F",
		X"51",X"20",X"12",X"20",X"31",X"0F",X"61",X"10",X"12",X"20",X"31",X"00",X"51",X"20",X"12",X"10",
		X"41",X"0F",X"51",X"20",X"12",X"20",X"31",X"0F",X"61",X"10",X"22",X"10",X"31",X"0F",X"61",X"20",
		X"12",X"20",X"31",X"0F",X"61",X"20",X"22",X"10",X"31",X"00",X"61",X"10",X"22",X"20",X"31",X"0F",
		X"61",X"20",X"12",X"20",X"31",X"0F",X"61",X"20",X"22",X"10",X"41",X"0F",X"71",X"10",X"22",X"20",
		X"31",X"0F",X"71",X"20",X"22",X"10",X"41",X"00",X"61",X"20",X"22",X"20",X"31",X"0F",X"61",X"20",
		X"22",X"20",X"41",X"0F",X"71",X"10",X"32",X"10",X"41",X"0F",X"71",X"20",X"22",X"20",X"41",X"0F",
		X"81",X"10",X"22",X"20",X"41",X"00",X"71",X"20",X"22",X"10",X"41",X"0F",X"81",X"10",X"22",X"20",
		X"41",X"0F",X"91",X"10",X"22",X"10",X"41",X"0F",X"91",X"20",X"12",X"20",X"41",X"10",X"12",X"00",
		X"91",X"10",X"12",X"20",X"41",X"0F",X"A1",X"10",X"12",X"10",X"51",X"0F",X"A1",X"40",X"41",X"0F",
		X"B1",X"10",X"12",X"10",X"51",X"10",X"12",X"0F",X"C1",X"30",X"41",X"0F",X"D1",X"20",X"51",X"00",
		X"C1",X"20",X"51",X"0F",X"D1",X"20",X"41",X"0F",X"E1",X"10",X"51",X"10",X"12",X"0F",X"F1",X"51",
		X"00",X"81",X"10",X"B1",X"10",X"12",X"0F",X"81",X"20",X"A1",X"0F",X"91",X"20",X"A1",X"10",X"12",
		X"0F",X"91",X"30",X"91",X"0F",X"91",X"30",X"A1",X"10",X"12",X"00",X"91",X"10",X"12",X"10",X"91",
		X"0F",X"91",X"20",X"12",X"10",X"91",X"10",X"12",X"0F",X"91",X"20",X"12",X"20",X"81",X"0F",X"91",
		X"20",X"22",X"10",X"91",X"10",X"12",X"0F",X"A1",X"10",X"32",X"10",X"81",X"00",X"91",X"20",X"32",
		X"10",X"81",X"10",X"12",X"0F",X"91",X"20",X"32",X"20",X"71",X"0F",X"A1",X"10",X"42",X"10",X"81",
		X"10",X"12",X"0F",X"A1",X"20",X"42",X"10",X"71",X"0F",X"A1",X"20",X"42",X"20",X"61",X"20",X"12",
		X"00",X"A1",X"10",X"52",X"10",X"71",X"10",X"12",X"0F",X"A1",X"20",X"42",X"20",X"61",X"20",X"12",
		X"0F",X"A1",X"20",X"52",X"10",X"71",X"10",X"12",X"0F",X"B1",X"10",X"52",X"20",X"61",X"20",X"12",
		X"0F",X"B1",X"20",X"42",X"20",X"71",X"10",X"12",X"00",X"A1",X"20",X"52",X"10",X"71",X"20",X"12",
		X"0F",X"B1",X"10",X"52",X"20",X"61",X"20",X"12",X"0F",X"B1",X"20",X"42",X"20",X"71",X"10",X"22",
		X"0F",X"B1",X"20",X"52",X"10",X"71",X"20",X"12",X"0F",X"B1",X"20",X"52",X"20",X"71",X"10",X"22",
		X"00",X"B1",X"10",X"52",X"20",X"71",X"20",X"12",X"0F",X"B1",X"20",X"52",X"10",X"81",X"10",X"22",
		X"0F",X"B1",X"20",X"52",X"20",X"71",X"20",X"12",X"0F",X"B1",X"20",X"52",X"20",X"71",X"20",X"22",
		X"0F",X"C1",X"10",X"62",X"10",X"81",X"10",X"22",X"00",X"B1",X"20",X"52",X"20",X"71",X"20",X"22",
		X"0F",X"B1",X"20",X"52",X"20",X"81",X"10",X"22",X"0F",X"B1",X"20",X"62",X"10",X"81",X"20",X"22",
		X"0F",X"C1",X"10",X"62",X"20",X"81",X"10",X"22",X"0F",X"C1",X"20",X"52",X"20",X"81",X"20",X"22",
		X"00",X"B1",X"20",X"62",X"10",X"91",X"10",X"22",X"0F",X"C1",X"10",X"62",X"20",X"81",X"20",X"22",
		X"0F",X"C1",X"20",X"62",X"10",X"91",X"10",X"22",X"0F",X"C1",X"20",X"62",X"20",X"81",X"20",X"22",
		X"0F",X"D1",X"10",X"72",X"10",X"81",X"20",X"22",X"00",X"C1",X"20",X"62",X"20",X"81",X"10",X"32",
		X"0F",X"C1",X"20",X"62",X"20",X"81",X"20",X"22",X"0F",X"D1",X"10",X"72",X"10",X"91",X"10",X"32",
		X"0F",X"D1",X"20",X"62",X"20",X"81",X"20",X"22",X"0F",X"D1",X"20",X"72",X"10",X"91",X"10",X"32",
		X"00",X"E0",X"82",X"B0",X"32",X"00",X"D2",X"10",X"82",X"10",X"92",X"10",X"32",X"00",X"D2",X"10",
		X"82",X"10",X"92",X"10",X"32",X"00",X"D2",X"10",X"82",X"10",X"92",X"10",X"32",X"00",X"D2",X"10",
		X"82",X"10",X"92",X"10",X"32",X"00",X"D2",X"10",X"82",X"10",X"92",X"10",X"32",X"00",X"D2",X"10",
		X"82",X"10",X"92",X"10",X"32",X"00",X"D2",X"10",X"72",X"20",X"92",X"10",X"32",X"00",X"D2",X"10",
		X"72",X"20",X"92",X"10",X"32",X"00",X"D2",X"10",X"62",X"30",X"92",X"10",X"32",X"00",X"D2",X"10",
		X"62",X"30",X"92",X"10",X"32",X"00",X"D2",X"10",X"52",X"40",X"92",X"10",X"32",X"00",X"D2",X"10",
		X"52",X"40",X"92",X"10",X"32",X"00",X"D2",X"10",X"42",X"50",X"92",X"10",X"32",X"00",X"D2",X"10",
		X"42",X"50",X"92",X"10",X"22",X"00",X"D2",X"10",X"32",X"60",X"92",X"10",X"22",X"00",X"D2",X"10",
		X"32",X"60",X"92",X"10",X"22",X"00",X"D2",X"10",X"22",X"70",X"92",X"10",X"12",X"00",X"D2",X"10",
		X"22",X"70",X"92",X"10",X"12",X"00",X"D2",X"10",X"12",X"80",X"92",X"10",X"12",X"00",X"D2",X"10",
		X"12",X"80",X"92",X"FF",X"B1",X"0F",X"C1",X"00",X"B1",X"0F",X"C1",X"00",X"C1",X"0F",X"61",X"00",
		X"51",X"20",X"62",X"0F",X"61",X"20",X"62",X"00",X"61",X"20",X"62",X"0F",X"61",X"30",X"62",X"00",
		X"61",X"10",X"12",X"10",X"62",X"0F",X"61",X"20",X"12",X"00",X"61",X"10",X"22",X"0F",X"71",X"10",
		X"22",X"00",X"61",X"20",X"22",X"0F",X"71",X"10",X"22",X"00",X"71",X"10",X"22",X"0F",X"71",X"20",
		X"22",X"00",X"71",X"10",X"22",X"0F",X"71",X"20",X"22",X"00",X"71",X"10",X"32",X"0F",X"71",X"20",
		X"22",X"00",X"71",X"10",X"32",X"0F",X"71",X"20",X"32",X"00",X"71",X"10",X"32",X"0F",X"71",X"20",
		X"32",X"00",X"71",X"10",X"42",X"0F",X"81",X"10",X"32",X"00",X"71",X"20",X"32",X"0F",X"81",X"10",
		X"42",X"00",X"71",X"20",X"32",X"0F",X"81",X"10",X"42",X"00",X"81",X"10",X"42",X"0F",X"81",X"20",
		X"32",X"00",X"81",X"0F",X"F1",X"31",X"00",X"F1",X"21",X"0F",X"F1",X"31",X"10",X"12",X"0F",X"F1",
		X"41",X"10",X"12",X"00",X"F1",X"31",X"20",X"12",X"0F",X"F1",X"41",X"10",X"22",X"00",X"F1",X"41",
		X"10",X"22",X"0F",X"F1",X"41",X"20",X"22",X"00",X"F1",X"41",X"10",X"32",X"0F",X"A1",X"B0",X"32",
		X"00",X"91",X"20",X"92",X"10",X"32",X"0F",X"A1",X"10",X"A2",X"10",X"32",X"00",X"91",X"20",X"A2",
		X"10",X"32",X"0F",X"A1",X"20",X"A2",X"10",X"22",X"00",X"A1",X"20",X"A2",X"10",X"22",X"0F",X"A1",
		X"30",X"A2",X"10",X"22",X"00",X"A1",X"10",X"12",X"10",X"A2",X"10",X"12",X"0F",X"B1",X"10",X"12",
		X"10",X"A2",X"10",X"12",X"00",X"A1",X"20",X"12",X"10",X"A2",X"10",X"12",X"0F",X"B1",X"10",X"22",
		X"10",X"A2",X"00",X"A1",X"20",X"22",X"10",X"A2",X"0F",X"B1",X"10",X"32",X"00",X"B1",X"10",X"32",
		X"0F",X"B1",X"20",X"32",X"00",X"B1",X"10",X"42",X"0F",X"B1",X"20",X"32",X"00",X"B1",X"10",X"42",
		X"0F",X"B1",X"20",X"42",X"00",X"B1",X"10",X"52",X"0F",X"C1",X"10",X"42",X"00",X"B1",X"20",X"42",
		X"0F",X"C1",X"10",X"52",X"00",X"B1",X"20",X"42",X"0F",X"C1",X"10",X"52",X"00",X"B1",X"20",X"52",
		X"0F",X"C1",X"10",X"52",X"00",X"C1",X"10",X"52",X"0F",X"C1",X"20",X"52",X"00",X"C1",X"10",X"52",
		X"0F",X"C1",X"20",X"52",X"00",X"C1",X"10",X"62",X"0F",X"C1",X"20",X"52",X"00",X"C1",X"10",X"62",
		X"0F",X"D1",X"10",X"62",X"00",X"C1",X"20",X"52",X"0F",X"D1",X"10",X"62",X"00",X"D1",X"10",X"62",
		X"0F",X"D1",X"20",X"62",X"00",X"D1",X"10",X"62",X"0F",X"D1",X"20",X"62",X"00",X"D1",X"10",X"72",
		X"0F",X"E1",X"10",X"62",X"00",X"F0",X"62",X"00",X"E2",X"10",X"62",X"00",X"E2",X"10",X"52",X"00",
		X"E2",X"10",X"52",X"00",X"E2",X"10",X"52",X"00",X"E2",X"10",X"42",X"00",X"E2",X"10",X"42",X"00",
		X"E2",X"10",X"42",X"00",X"E2",X"10",X"42",X"00",X"E2",X"10",X"32",X"00",X"E2",X"10",X"32",X"00",
		X"E2",X"10",X"32",X"00",X"E2",X"10",X"22",X"00",X"E2",X"10",X"22",X"00",X"E2",X"10",X"22",X"00",
		X"E2",X"10",X"12",X"00",X"E2",X"10",X"12",X"00",X"E2",X"10",X"12",X"00",X"E2",X"10",X"12",X"00",
		X"E2",X"00",X"E2",X"FF",X"B1",X"00",X"B1",X"00",X"B1",X"00",X"B1",X"0F",X"C1",X"00",X"51",X"00",
		X"51",X"10",X"62",X"00",X"51",X"10",X"62",X"0F",X"51",X"20",X"62",X"00",X"51",X"20",X"62",X"00",
		X"51",X"20",X"62",X"00",X"51",X"0F",X"61",X"10",X"12",X"00",X"61",X"10",X"12",X"00",X"61",X"10",
		X"12",X"00",X"61",X"10",X"12",X"00",X"61",X"10",X"12",X"0F",X"61",X"20",X"12",X"00",X"61",X"10",
		X"22",X"00",X"61",X"10",X"12",X"00",X"61",X"10",X"12",X"0F",X"71",X"10",X"12",X"00",X"71",X"10",
		X"12",X"00",X"71",X"10",X"12",X"00",X"71",X"10",X"12",X"00",X"71",X"10",X"12",X"0F",X"81",X"10",
		X"12",X"00",X"71",X"20",X"12",X"00",X"71",X"10",X"22",X"00",X"71",X"10",X"12",X"0F",X"81",X"10",
		X"12",X"00",X"81",X"10",X"12",X"00",X"81",X"10",X"12",X"00",X"81",X"10",X"12",X"00",X"81",X"0F",
		X"F1",X"31",X"00",X"F1",X"31",X"00",X"F1",X"31",X"10",X"12",X"00",X"F1",X"31",X"10",X"12",X"00",
		X"F1",X"31",X"10",X"12",X"0F",X"F1",X"41",X"10",X"12",X"00",X"F1",X"41",X"10",X"12",X"00",X"F1",
		X"41",X"10",X"12",X"00",X"F1",X"41",X"10",X"12",X"0F",X"F1",X"51",X"10",X"12",X"00",X"91",X"C0",
		X"12",X"00",X"91",X"10",X"A2",X"10",X"12",X"00",X"91",X"10",X"A2",X"10",X"12",X"00",X"91",X"10",
		X"A2",X"10",X"12",X"0F",X"A1",X"10",X"A2",X"10",X"12",X"00",X"A1",X"10",X"A2",X"10",X"12",X"00",
		X"A1",X"10",X"A2",X"10",X"12",X"00",X"A1",X"10",X"A2",X"10",X"12",X"0F",X"B1",X"10",X"A2",X"10",
		X"12",X"00",X"B1",X"10",X"A2",X"10",X"12",X"00",X"A1",X"20",X"A2",X"00",X"A1",X"0F",X"B1",X"10",
		X"12",X"00",X"B1",X"10",X"12",X"00",X"B1",X"10",X"12",X"00",X"B1",X"10",X"12",X"0F",X"C1",X"10",
		X"12",X"00",X"C1",X"10",X"12",X"00",X"C1",X"10",X"12",X"00",X"C1",X"10",X"12",X"00",X"B1",X"20",
		X"12",X"0F",X"C1",X"10",X"22",X"00",X"C1",X"10",X"12",X"00",X"C1",X"10",X"12",X"00",X"C1",X"10",
		X"12",X"00",X"C1",X"10",X"12",X"0F",X"D1",X"10",X"12",X"00",X"D1",X"10",X"12",X"00",X"D1",X"00",
		X"F1",X"F1",X"0F",X"F1",X"F1",X"11",X"00",X"F1",X"F1",X"11",X"00",X"F1",X"F1",X"11",X"00",X"F1",
		X"F1",X"11",X"0F",X"F1",X"F1",X"21",X"00",X"F1",X"F1",X"31",X"00",X"F1",X"F1",X"31",X"00",X"F1",
		X"F1",X"31",X"0F",X"F1",X"F1",X"41",X"00",X"F1",X"F1",X"41",X"00",X"F1",X"F1",X"41",X"0F",X"F1",
		X"F1",X"51",X"00",X"00",X"F2",X"F2",X"52",X"00",X"F2",X"F2",X"52",X"00",X"F2",X"F2",X"52",X"00",
		X"F2",X"F2",X"52",X"00",X"F2",X"F2",X"52",X"00",X"F2",X"F2",X"52",X"00",X"F2",X"F2",X"52",X"00",
		X"F2",X"F2",X"52",X"00",X"F2",X"F2",X"52",X"00",X"F2",X"F2",X"52",X"00",X"F2",X"F2",X"52",X"00",
		X"F2",X"F2",X"52",X"00",X"F2",X"F2",X"52",X"00",X"F2",X"F2",X"52",X"00",X"F2",X"F2",X"52",X"00",
		X"F2",X"F2",X"52",X"00",X"F2",X"F2",X"52",X"00",X"F2",X"F2",X"52",X"00",X"F2",X"F2",X"52",X"00",
		X"F2",X"F2",X"52",X"FF",X"91",X"00",X"A1",X"00",X"B1",X"00",X"C1",X"00",X"C1",X"00",X"51",X"40",
		X"31",X"00",X"51",X"10",X"22",X"10",X"31",X"01",X"41",X"20",X"12",X"20",X"31",X"0E",X"12",X"10",
		X"51",X"10",X"22",X"10",X"31",X"00",X"12",X"10",X"51",X"10",X"22",X"10",X"31",X"00",X"12",X"10",
		X"51",X"10",X"22",X"10",X"41",X"00",X"12",X"10",X"51",X"20",X"12",X"20",X"31",X"00",X"12",X"10",
		X"51",X"20",X"22",X"10",X"31",X"00",X"12",X"10",X"51",X"20",X"22",X"10",X"41",X"00",X"12",X"10",
		X"61",X"20",X"12",X"10",X"41",X"00",X"12",X"10",X"61",X"20",X"12",X"20",X"31",X"00",X"12",X"20",
		X"51",X"20",X"22",X"10",X"41",X"00",X"22",X"10",X"51",X"20",X"22",X"10",X"41",X"01",X"12",X"10",
		X"51",X"30",X"12",X"10",X"41",X"00",X"12",X"10",X"61",X"20",X"12",X"20",X"41",X"00",X"12",X"10",
		X"61",X"20",X"22",X"10",X"41",X"00",X"12",X"10",X"61",X"20",X"22",X"10",X"41",X"00",X"12",X"10",
		X"61",X"20",X"22",X"10",X"51",X"00",X"12",X"10",X"71",X"20",X"12",X"20",X"41",X"00",X"12",X"10",
		X"71",X"20",X"22",X"10",X"41",X"00",X"12",X"10",X"71",X"20",X"22",X"10",X"51",X"00",X"12",X"10",
		X"71",X"20",X"22",X"20",X"41",X"00",X"12",X"20",X"61",X"20",X"32",X"10",X"51",X"00",X"22",X"10",
		X"71",X"20",X"22",X"10",X"51",X"01",X"12",X"10",X"71",X"20",X"22",X"10",X"51",X"00",X"12",X"10",
		X"71",X"20",X"22",X"10",X"61",X"00",X"12",X"10",X"71",X"20",X"22",X"10",X"61",X"00",X"12",X"10",
		X"81",X"10",X"12",X"20",X"61",X"00",X"12",X"10",X"81",X"30",X"71",X"00",X"12",X"10",X"81",X"20",
		X"81",X"00",X"12",X"10",X"F1",X"31",X"00",X"12",X"10",X"F1",X"31",X"00",X"12",X"10",X"F1",X"21",
		X"00",X"12",X"10",X"F1",X"21",X"00",X"12",X"10",X"F1",X"11",X"00",X"12",X"10",X"F1",X"00",X"12",
		X"20",X"F1",X"11",X"00",X"22",X"10",X"F1",X"21",X"01",X"12",X"10",X"F1",X"31",X"00",X"12",X"10",
		X"F1",X"41",X"00",X"12",X"10",X"91",X"20",X"91",X"00",X"12",X"10",X"91",X"30",X"91",X"00",X"12",
		X"10",X"91",X"10",X"12",X"20",X"91",X"00",X"12",X"10",X"91",X"20",X"12",X"20",X"81",X"00",X"12",
		X"10",X"A1",X"10",X"22",X"20",X"81",X"00",X"12",X"10",X"A1",X"10",X"32",X"20",X"71",X"00",X"12",
		X"10",X"A1",X"10",X"42",X"10",X"81",X"00",X"12",X"10",X"A1",X"10",X"42",X"20",X"71",X"00",X"12",
		X"10",X"A1",X"20",X"42",X"10",X"81",X"00",X"12",X"20",X"A1",X"10",X"42",X"20",X"71",X"00",X"22",
		X"10",X"A1",X"10",X"52",X"10",X"71",X"01",X"12",X"10",X"A1",X"20",X"42",X"10",X"81",X"00",X"12",
		X"10",X"A1",X"20",X"42",X"20",X"71",X"00",X"12",X"10",X"A1",X"20",X"52",X"10",X"71",X"00",X"12",
		X"10",X"A1",X"30",X"42",X"10",X"81",X"00",X"12",X"10",X"B1",X"20",X"42",X"20",X"71",X"00",X"12",
		X"10",X"B1",X"20",X"52",X"10",X"81",X"00",X"12",X"10",X"B1",X"20",X"52",X"10",X"81",X"00",X"12",
		X"10",X"B1",X"30",X"42",X"10",X"81",X"00",X"12",X"10",X"B1",X"30",X"42",X"20",X"81",X"00",X"12",
		X"10",X"C1",X"20",X"42",X"20",X"81",X"00",X"12",X"10",X"C1",X"20",X"52",X"10",X"81",X"00",X"12",
		X"20",X"B1",X"30",X"42",X"20",X"81",X"00",X"22",X"10",X"B1",X"30",X"52",X"10",X"81",X"01",X"12",
		X"10",X"B1",X"30",X"52",X"10",X"91",X"00",X"12",X"10",X"C1",X"20",X"52",X"20",X"81",X"00",X"12",
		X"10",X"C1",X"30",X"52",X"10",X"81",X"00",X"12",X"10",X"C1",X"30",X"52",X"10",X"91",X"00",X"12",
		X"10",X"C1",X"30",X"52",X"10",X"91",X"00",X"12",X"10",X"D1",X"20",X"52",X"20",X"81",X"00",X"12",
		X"10",X"D1",X"30",X"52",X"10",X"91",X"00",X"12",X"10",X"D1",X"30",X"52",X"10",X"91",X"00",X"12",
		X"10",X"D1",X"30",X"52",X"10",X"91",X"00",X"12",X"10",X"E1",X"20",X"52",X"20",X"91",X"00",X"12",
		X"10",X"E1",X"30",X"52",X"10",X"91",X"00",X"12",X"20",X"D1",X"30",X"52",X"10",X"91",X"00",X"22",
		X"10",X"D1",X"30",X"52",X"10",X"A1",X"01",X"12",X"10",X"E1",X"20",X"52",X"20",X"91",X"00",X"12",
		X"10",X"E1",X"30",X"52",X"10",X"91",X"00",X"12",X"10",X"E1",X"30",X"52",X"10",X"A1",X"00",X"12",
		X"10",X"E1",X"30",X"52",X"20",X"91",X"00",X"12",X"10",X"F1",X"20",X"62",X"10",X"A1",X"00",X"12",
		X"F0",X"40",X"52",X"00",X"12",X"10",X"F2",X"30",X"52",X"10",X"A2",X"00",X"12",X"10",X"F2",X"30",
		X"52",X"10",X"A2",X"00",X"12",X"10",X"F2",X"30",X"52",X"10",X"A2",X"00",X"12",X"10",X"F2",X"40",
		X"42",X"10",X"A2",X"00",X"12",X"10",X"F2",X"40",X"42",X"10",X"A2",X"00",X"12",X"10",X"F2",X"40",
		X"42",X"10",X"A2",X"00",X"12",X"10",X"F2",X"40",X"42",X"10",X"A2",X"00",X"12",X"10",X"F2",X"50",
		X"32",X"10",X"A2",X"00",X"12",X"10",X"F2",X"50",X"32",X"10",X"A2",X"00",X"12",X"10",X"F2",X"50",
		X"32",X"10",X"A2",X"00",X"12",X"10",X"F2",X"50",X"32",X"10",X"A2",X"00",X"12",X"10",X"F2",X"60",
		X"22",X"10",X"A2",X"00",X"12",X"10",X"F2",X"60",X"22",X"10",X"A2",X"02",X"F2",X"60",X"22",X"10",
		X"A2",X"00",X"F2",X"60",X"22",X"10",X"A2",X"00",X"F2",X"70",X"12",X"10",X"A2",X"00",X"F2",X"70",
		X"12",X"10",X"A2",X"00",X"F2",X"70",X"12",X"10",X"A2",X"00",X"F2",X"70",X"12",X"10",X"A2",X"00",
		X"F2",X"90",X"A2",X"FF",X"41",X"30",X"31",X"01",X"31",X"40",X"21",X"00",X"41",X"20",X"12",X"10",
		X"21",X"01",X"31",X"20",X"12",X"10",X"21",X"0E",X"12",X"10",X"41",X"10",X"12",X"20",X"21",X"00",
		X"12",X"20",X"31",X"20",X"12",X"10",X"31",X"01",X"12",X"10",X"41",X"10",X"12",X"20",X"21",X"00",
		X"12",X"10",X"41",X"10",X"22",X"10",X"31",X"00",X"12",X"20",X"31",X"20",X"12",X"20",X"31",X"01",
		X"12",X"10",X"41",X"10",X"22",X"20",X"21",X"00",X"12",X"10",X"41",X"20",X"22",X"10",X"31",X"00",
		X"12",X"20",X"41",X"10",X"22",X"20",X"31",X"01",X"12",X"10",X"41",X"20",X"22",X"10",X"31",X"00",
		X"12",X"10",X"51",X"10",X"22",X"20",X"31",X"00",X"12",X"20",X"41",X"20",X"22",X"20",X"31",X"01",
		X"12",X"10",X"51",X"10",X"32",X"10",X"31",X"00",X"12",X"10",X"51",X"20",X"22",X"20",X"31",X"00",
		X"12",X"20",X"51",X"10",X"32",X"10",X"41",X"01",X"12",X"10",X"51",X"20",X"22",X"20",X"31",X"00",
		X"12",X"10",X"61",X"10",X"32",X"10",X"41",X"00",X"12",X"20",X"51",X"20",X"22",X"20",X"41",X"01",
		X"12",X"10",X"61",X"10",X"32",X"10",X"41",X"00",X"12",X"10",X"61",X"20",X"22",X"20",X"41",X"00",
		X"12",X"20",X"61",X"10",X"32",X"10",X"51",X"01",X"12",X"10",X"61",X"20",X"22",X"20",X"41",X"00",
		X"12",X"20",X"61",X"10",X"32",X"10",X"51",X"01",X"12",X"10",X"61",X"20",X"22",X"20",X"51",X"00",
		X"12",X"10",X"71",X"20",X"22",X"10",X"51",X"00",X"12",X"20",X"71",X"20",X"12",X"20",X"51",X"01",
		X"12",X"10",X"81",X"20",X"12",X"20",X"51",X"00",X"12",X"10",X"91",X"20",X"12",X"10",X"51",X"00",
		X"12",X"20",X"91",X"40",X"51",X"00",X"22",X"10",X"A1",X"30",X"51",X"00",X"22",X"10",X"C1",X"20",
		X"51",X"00",X"22",X"20",X"C1",X"20",X"51",X"00",X"32",X"10",X"D1",X"10",X"51",X"00",X"32",X"20",
		X"D1",X"10",X"51",X"00",X"42",X"10",X"F1",X"51",X"00",X"42",X"10",X"F1",X"51",X"00",X"42",X"20",
		X"F1",X"51",X"00",X"52",X"10",X"F1",X"61",X"00",X"52",X"10",X"91",X"10",X"B1",X"01",X"42",X"20",
		X"91",X"10",X"B1",X"01",X"42",X"10",X"91",X"20",X"B1",X"01",X"32",X"10",X"A1",X"20",X"A1",X"01",
		X"22",X"20",X"91",X"30",X"A1",X"01",X"22",X"10",X"A1",X"10",X"12",X"10",X"A1",X"00",X"22",X"10",
		X"A1",X"40",X"91",X"01",X"12",X"20",X"A1",X"10",X"12",X"20",X"91",X"00",X"22",X"10",X"A1",X"20",
		X"12",X"20",X"91",X"01",X"12",X"20",X"A1",X"10",X"22",X"10",X"91",X"00",X"22",X"10",X"A1",X"20",
		X"12",X"20",X"91",X"01",X"12",X"10",X"B1",X"10",X"22",X"20",X"81",X"00",X"12",X"20",X"A1",X"20",
		X"22",X"20",X"81",X"00",X"22",X"10",X"B1",X"10",X"32",X"20",X"81",X"01",X"12",X"20",X"A1",X"20",
		X"32",X"20",X"71",X"00",X"22",X"10",X"B1",X"10",X"42",X"20",X"71",X"00",X"22",X"20",X"A1",X"20",
		X"42",X"20",X"71",X"01",X"22",X"10",X"B1",X"10",X"52",X"20",X"61",X"00",X"22",X"10",X"B1",X"20",
		X"42",X"20",X"71",X"01",X"12",X"20",X"B1",X"10",X"42",X"30",X"71",X"00",X"22",X"10",X"B1",X"20",
		X"32",X"10",X"12",X"10",X"71",X"00",X"22",X"10",X"C1",X"10",X"32",X"10",X"12",X"20",X"71",X"01",
		X"12",X"20",X"B1",X"20",X"22",X"10",X"22",X"10",X"81",X"00",X"22",X"10",X"C1",X"10",X"22",X"10",
		X"22",X"20",X"71",X"00",X"22",X"20",X"B1",X"20",X"12",X"10",X"32",X"10",X"81",X"01",X"22",X"10",
		X"C1",X"10",X"12",X"10",X"32",X"20",X"81",X"00",X"22",X"10",X"C1",X"30",X"42",X"10",X"81",X"01",
		X"12",X"20",X"C1",X"20",X"42",X"20",X"81",X"00",X"22",X"10",X"C1",X"20",X"52",X"10",X"91",X"00",
		X"22",X"20",X"C1",X"10",X"52",X"20",X"81",X"01",X"22",X"10",X"C1",X"20",X"52",X"20",X"81",X"00",
		X"22",X"10",X"D1",X"10",X"62",X"10",X"91",X"00",X"22",X"20",X"C1",X"20",X"52",X"20",X"81",X"01",
		X"22",X"10",X"D1",X"10",X"62",X"10",X"91",X"00",X"22",X"20",X"C1",X"20",X"52",X"20",X"91",X"00",
		X"32",X"10",X"D1",X"10",X"62",X"10",X"91",X"01",X"22",X"10",X"D1",X"20",X"52",X"20",X"91",X"00",
		X"22",X"20",X"D1",X"10",X"62",X"10",X"A1",X"00",X"32",X"10",X"D1",X"20",X"52",X"20",X"91",X"01",
		X"22",X"10",X"E1",X"10",X"62",X"10",X"A1",X"00",X"22",X"20",X"D1",X"20",X"52",X"20",X"A1",X"00",
		X"32",X"10",X"E1",X"10",X"62",X"10",X"A1",X"01",X"22",X"20",X"D1",X"20",X"52",X"20",X"A1",X"00",
		X"32",X"10",X"E1",X"10",X"62",X"10",X"B1",X"01",X"22",X"20",X"D1",X"20",X"52",X"20",X"A1",X"00",
		X"32",X"10",X"E1",X"10",X"62",X"10",X"B1",X"00",X"32",X"F0",X"10",X"62",X"00",X"32",X"10",X"E2",
		X"10",X"62",X"10",X"B2",X"00",X"32",X"10",X"E2",X"10",X"62",X"10",X"B2",X"00",X"32",X"10",X"E2",
		X"10",X"62",X"10",X"B2",X"00",X"32",X"10",X"E2",X"10",X"62",X"10",X"B2",X"00",X"32",X"10",X"E2",
		X"10",X"62",X"10",X"B2",X"00",X"32",X"10",X"E2",X"10",X"62",X"10",X"B2",X"00",X"32",X"10",X"E2",
		X"10",X"62",X"10",X"B2",X"00",X"32",X"10",X"E2",X"10",X"62",X"10",X"B2",X"00",X"32",X"10",X"E2",
		X"10",X"62",X"10",X"B2",X"00",X"32",X"10",X"E2",X"20",X"52",X"10",X"B2",X"00",X"32",X"10",X"E2",
		X"20",X"52",X"10",X"B2",X"00",X"32",X"10",X"E2",X"30",X"42",X"10",X"B2",X"00",X"32",X"10",X"E2",
		X"30",X"42",X"10",X"B2",X"01",X"22",X"10",X"E2",X"40",X"32",X"10",X"B2",X"00",X"22",X"10",X"E2",
		X"40",X"32",X"10",X"B2",X"00",X"22",X"10",X"E2",X"50",X"22",X"10",X"B2",X"01",X"12",X"10",X"E2",
		X"50",X"22",X"10",X"B2",X"00",X"12",X"10",X"E2",X"60",X"12",X"10",X"B2",X"00",X"12",X"10",X"E2",
		X"60",X"12",X"10",X"B2",X"02",X"E2",X"80",X"B2",X"FF",X"31",X"0F",X"71",X"0F",X"A1",X"00",X"B1",
		X"00",X"41",X"40",X"41",X"00",X"41",X"50",X"41",X"01",X"41",X"50",X"41",X"00",X"51",X"20",X"12",
		X"20",X"41",X"01",X"51",X"20",X"12",X"20",X"41",X"01",X"51",X"10",X"22",X"20",X"41",X"00",X"51",
		X"20",X"22",X"20",X"41",X"01",X"51",X"20",X"22",X"20",X"41",X"01",X"51",X"20",X"22",X"10",X"51",
		X"01",X"51",X"20",X"12",X"20",X"51",X"0E",X"12",X"10",X"61",X"10",X"22",X"20",X"51",X"03",X"51",
		X"20",X"22",X"20",X"51",X"01",X"51",X"20",X"22",X"20",X"51",X"0E",X"12",X"10",X"61",X"20",X"22",
		X"20",X"51",X"03",X"61",X"20",X"22",X"20",X"51",X"01",X"61",X"10",X"32",X"10",X"61",X"0E",X"12",
		X"10",X"61",X"20",X"22",X"20",X"61",X"03",X"61",X"20",X"22",X"20",X"61",X"01",X"61",X"20",X"22",
		X"20",X"61",X"0E",X"12",X"20",X"61",X"20",X"22",X"20",X"61",X"01",X"12",X"10",X"71",X"10",X"32",
		X"20",X"61",X"01",X"20",X"61",X"20",X"32",X"20",X"61",X"00",X"12",X"20",X"61",X"20",X"32",X"10",
		X"71",X"01",X"12",X"10",X"71",X"20",X"22",X"20",X"71",X"01",X"20",X"71",X"20",X"22",X"20",X"71",
		X"00",X"12",X"10",X"81",X"10",X"32",X"20",X"71",X"01",X"20",X"71",X"20",X"32",X"20",X"71",X"00",
		X"12",X"20",X"71",X"20",X"32",X"20",X"71",X"01",X"12",X"20",X"71",X"20",X"32",X"20",X"71",X"01",
		X"12",X"10",X"81",X"20",X"32",X"20",X"71",X"00",X"12",X"20",X"81",X"20",X"32",X"20",X"71",X"01",
		X"12",X"20",X"81",X"10",X"42",X"20",X"71",X"01",X"12",X"10",X"81",X"20",X"42",X"20",X"71",X"00",
		X"12",X"20",X"81",X"20",X"42",X"10",X"81",X"01",X"12",X"20",X"81",X"20",X"32",X"20",X"81",X"01",
		X"12",X"10",X"91",X"20",X"32",X"20",X"81",X"00",X"12",X"20",X"91",X"20",X"32",X"20",X"81",X"01",
		X"12",X"20",X"91",X"10",X"42",X"20",X"81",X"01",X"12",X"20",X"81",X"20",X"42",X"20",X"81",X"00",
		X"22",X"10",X"91",X"20",X"42",X"20",X"81",X"01",X"12",X"20",X"91",X"20",X"42",X"20",X"81",X"01",
		X"12",X"20",X"91",X"20",X"42",X"20",X"81",X"00",X"22",X"10",X"A1",X"10",X"52",X"20",X"81",X"01",
		X"12",X"20",X"91",X"20",X"52",X"20",X"81",X"01",X"12",X"10",X"A1",X"20",X"52",X"20",X"81",X"00",
		X"12",X"20",X"A1",X"20",X"52",X"20",X"81",X"01",X"12",X"20",X"A1",X"10",X"62",X"20",X"81",X"00",
		X"22",X"20",X"91",X"20",X"62",X"20",X"81",X"01",X"22",X"10",X"A1",X"20",X"62",X"20",X"81",X"01",
		X"12",X"20",X"A1",X"20",X"62",X"10",X"91",X"00",X"22",X"20",X"A1",X"20",X"52",X"20",X"91",X"01",
		X"22",X"10",X"B1",X"10",X"62",X"20",X"91",X"01",X"12",X"20",X"A1",X"20",X"62",X"20",X"91",X"00",
		X"22",X"20",X"A1",X"20",X"62",X"20",X"91",X"01",X"22",X"10",X"B1",X"20",X"62",X"20",X"91",X"01",
		X"12",X"20",X"B1",X"20",X"62",X"20",X"91",X"00",X"22",X"20",X"B1",X"20",X"62",X"20",X"91",X"01",
		X"22",X"10",X"C1",X"10",X"72",X"10",X"A1",X"01",X"12",X"20",X"B1",X"20",X"62",X"20",X"A1",X"00",
		X"22",X"20",X"B1",X"20",X"62",X"20",X"A1",X"01",X"22",X"20",X"B1",X"20",X"62",X"20",X"A1",X"01",
		X"22",X"20",X"B1",X"20",X"62",X"20",X"A1",X"00",X"32",X"10",X"C1",X"20",X"62",X"20",X"A1",X"01",
		X"22",X"20",X"C1",X"20",X"62",X"20",X"A1",X"01",X"22",X"20",X"C1",X"20",X"62",X"20",X"A1",X"00",
		X"32",X"10",X"D1",X"20",X"62",X"10",X"A1",X"01",X"22",X"20",X"D1",X"20",X"52",X"20",X"A1",X"01",
		X"22",X"20",X"D1",X"30",X"42",X"10",X"A1",X"00",X"32",X"10",X"F1",X"30",X"12",X"20",X"B1",X"01",
		X"22",X"20",X"F1",X"11",X"30",X"C1",X"01",X"22",X"20",X"F1",X"F1",X"00",X"32",X"20",X"F1",X"F1",
		X"01",X"32",X"20",X"F1",X"E1",X"01",X"32",X"20",X"F1",X"D1",X"00",X"42",X"20",X"F1",X"C1",X"01",
		X"42",X"20",X"F1",X"B1",X"01",X"42",X"20",X"F1",X"A1",X"00",X"52",X"20",X"F1",X"81",X"01",X"52",
		X"30",X"F1",X"61",X"10",X"12",X"01",X"62",X"30",X"F1",X"31",X"20",X"12",X"00",X"82",X"30",X"F1",
		X"11",X"10",X"22",X"01",X"92",X"30",X"D1",X"20",X"22",X"00",X"B2",X"30",X"A1",X"20",X"32",X"00",
		X"D2",X"C0",X"42",X"00",X"F2",X"E2",X"00",X"F2",X"E2",X"00",X"F2",X"E2",X"00",X"F2",X"E2",X"00",
		X"F2",X"E2",X"00",X"F2",X"E2",X"00",X"F2",X"E2",X"00",X"F2",X"E2",X"00",X"F2",X"E2",X"00",X"F2",
		X"D2",X"00",X"F2",X"D2",X"01",X"F2",X"C2",X"01",X"F2",X"B2",X"01",X"F2",X"92",X"01",X"F2",X"82",
		X"01",X"F2",X"72",X"01",X"F2",X"52",X"02",X"F2",X"22",X"02",X"E2",X"02",X"B2",X"FF",X"5F",X"34",
		X"56",X"A6",X"A0",X"81",X"FF",X"27",X"6D",X"85",X"F0",X"26",X"1A",X"48",X"48",X"48",X"48",X"47",
		X"47",X"47",X"47",X"6F",X"61",X"C6",X"01",X"AE",X"62",X"30",X"8B",X"AF",X"62",X"6A",X"E4",X"26",
		X"E0",X"1C",X"FE",X"35",X"D6",X"84",X"0F",X"C6",X"11",X"3D",X"A6",X"3F",X"44",X"44",X"44",X"44",
		X"5D",X"27",X"3A",X"34",X"16",X"1E",X"01",X"8B",X"14",X"46",X"1E",X"01",X"24",X"0F",X"C4",X"0F",
		X"EA",X"65",X"E7",X"84",X"E6",X"61",X"30",X"89",X"01",X"00",X"4A",X"27",X"19",X"81",X"02",X"25",
		X"0A",X"E7",X"84",X"30",X"89",X"01",X"00",X"80",X"02",X"20",X"F2",X"6F",X"65",X"4D",X"27",X"06",
		X"C4",X"F0",X"E7",X"84",X"E7",X"65",X"35",X"16",X"5F",X"30",X"8B",X"20",X"94",X"6F",X"61",X"5F",
		X"30",X"8B",X"20",X"8D",X"1A",X"01",X"35",X"D6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"49",X"4E",X"7E",X"49",X"96",X"7E",X"49",X"C1",X"7E",X"49",X"46",X"7E",X"49",X"8E",X"7E",
		X"49",X"B9",X"7E",X"4A",X"3F",X"7E",X"4A",X"2F",X"7E",X"4A",X"39",X"7E",X"4A",X"29",X"7E",X"49",
		X"D8",X"7E",X"49",X"24",X"34",X"76",X"8E",X"4A",X"94",X"1F",X"89",X"3A",X"3A",X"AE",X"84",X"4F",
		X"E6",X"84",X"C4",X"7F",X"BD",X"E0",X"5D",X"E6",X"80",X"2A",X"F5",X"44",X"40",X"8B",X"48",X"A7",
		X"62",X"35",X"76",X"7E",X"E0",X"10",X"34",X"67",X"10",X"8E",X"30",X"6A",X"20",X"06",X"34",X"67",
		X"10",X"8E",X"30",X"00",X"1A",X"FF",X"F7",X"C8",X"81",X"8D",X"02",X"35",X"E7",X"34",X"20",X"BF",
		X"C8",X"84",X"8C",X"90",X"00",X"22",X"1B",X"48",X"81",X"6A",X"25",X"02",X"86",X"5C",X"10",X"AE",
		X"A6",X"EC",X"A1",X"FD",X"C8",X"86",X"10",X"BF",X"C8",X"82",X"C6",X"1A",X"F7",X"C8",X"80",X"5F",
		X"30",X"8B",X"35",X"A0",X"84",X"0F",X"81",X"0A",X"2F",X"02",X"86",X"0A",X"20",X"CF",X"34",X"67",
		X"10",X"8E",X"30",X"6A",X"20",X"06",X"34",X"67",X"10",X"8E",X"30",X"00",X"1A",X"FF",X"F7",X"C8",
		X"81",X"CE",X"4A",X"94",X"1F",X"89",X"1E",X"31",X"3A",X"3A",X"1E",X"31",X"EE",X"C4",X"A6",X"C4",
		X"BD",X"49",X"5D",X"A6",X"C0",X"2A",X"F7",X"35",X"E7",X"34",X"67",X"10",X"8E",X"30",X"6A",X"20",
		X"06",X"34",X"67",X"10",X"8E",X"30",X"00",X"1A",X"FF",X"F7",X"C8",X"81",X"44",X"44",X"44",X"44",
		X"8D",X"B2",X"A6",X"61",X"8D",X"AE",X"35",X"E7",X"34",X"67",X"1F",X"23",X"10",X"8E",X"30",X"00",
		X"1A",X"FF",X"F7",X"C8",X"81",X"30",X"89",X"FD",X"00",X"5F",X"A6",X"C0",X"84",X"0F",X"8D",X"15",
		X"8D",X"11",X"8D",X"0F",X"8D",X"0D",X"5D",X"26",X"08",X"30",X"89",X"FD",X"00",X"4F",X"BD",X"49",
		X"84",X"35",X"E7",X"A6",X"C0",X"26",X"08",X"5D",X"26",X"05",X"30",X"89",X"06",X"00",X"39",X"5D",
		X"26",X"06",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"5C",X"34",X"06",X"44",X"44",X"44",X"44",X"BD",
		X"49",X"84",X"A6",X"E4",X"BD",X"49",X"84",X"35",X"86",X"34",X"66",X"C6",X"01",X"20",X"03",X"34",
		X"66",X"5F",X"E7",X"E4",X"CE",X"E0",X"25",X"20",X"0E",X"34",X"66",X"C6",X"01",X"20",X"03",X"34",
		X"66",X"5F",X"E7",X"E4",X"CE",X"E0",X"10",X"10",X"8E",X"58",X"7E",X"48",X"31",X"B6",X"EC",X"A1",
		X"27",X"02",X"AE",X"3E",X"EC",X"A1",X"6D",X"E4",X"27",X"01",X"5F",X"84",X"7F",X"AD",X"C4",X"6D",
		X"3E",X"2A",X"EB",X"35",X"04",X"35",X"E4",X"20",X"49",X"4E",X"46",X"45",X"52",X"4E",X"4F",X"20",
		X"2D",X"20",X"28",X"43",X"29",X"31",X"39",X"38",X"34",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",
		X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",
		X"4E",X"43",X"2E",X"20",X"52",X"47",X"52",X"57",X"52",X"6D",X"52",X"7B",X"52",X"85",X"52",X"8F",
		X"52",X"9F",X"52",X"B4",X"52",X"C7",X"52",X"CA",X"52",X"D2",X"52",X"E0",X"52",X"F7",X"53",X"13",
		X"53",X"2B",X"53",X"36",X"53",X"3D",X"53",X"44",X"53",X"4E",X"53",X"5E",X"53",X"67",X"53",X"72",
		X"53",X"7D",X"53",X"8D",X"58",X"13",X"58",X"1F",X"58",X"2A",X"58",X"38",X"58",X"45",X"58",X"51",
		X"53",X"9D",X"53",X"A7",X"53",X"BA",X"53",X"C9",X"53",X"DA",X"53",X"EA",X"53",X"F6",X"53",X"FE",
		X"54",X"13",X"54",X"23",X"54",X"36",X"4C",X"D1",X"54",X"47",X"54",X"5B",X"54",X"72",X"4C",X"DD",
		X"54",X"83",X"54",X"98",X"54",X"B2",X"54",X"C3",X"54",X"D2",X"54",X"E3",X"54",X"F3",X"55",X"0C",
		X"55",X"2B",X"55",X"47",X"55",X"59",X"55",X"72",X"55",X"8A",X"55",X"A2",X"55",X"B8",X"55",X"C2",
		X"55",X"DA",X"55",X"F0",X"56",X"04",X"56",X"21",X"56",X"24",X"56",X"2E",X"56",X"34",X"56",X"4D",
		X"56",X"55",X"56",X"6E",X"56",X"90",X"56",X"AB",X"56",X"B3",X"56",X"C9",X"56",X"D7",X"56",X"E5",
		X"56",X"ED",X"57",X"00",X"57",X"CC",X"57",X"DB",X"58",X"00",X"57",X"1E",X"57",X"35",X"57",X"48",
		X"57",X"55",X"57",X"65",X"57",X"98",X"57",X"BA",X"57",X"C3",X"58",X"5C",X"58",X"6A",X"58",X"77",
		X"52",X"40",X"52",X"3A",X"52",X"14",X"52",X"20",X"52",X"1C",X"51",X"FB",X"52",X"09",X"51",X"AD",
		X"51",X"B3",X"51",X"C0",X"51",X"C9",X"51",X"CB",X"51",X"E6",X"51",X"F0",X"51",X"89",X"51",X"94",
		X"51",X"A1",X"51",X"6B",X"51",X"75",X"51",X"7F",X"4D",X"8A",X"4D",X"9E",X"4D",X"B7",X"4D",X"DB",
		X"4D",X"F8",X"4E",X"0A",X"4E",X"2E",X"4E",X"50",X"4E",X"67",X"4E",X"82",X"4E",X"9B",X"4E",X"B5",
		X"4E",X"C8",X"4E",X"E3",X"4C",X"F2",X"4D",X"0E",X"4D",X"22",X"4F",X"0F",X"4F",X"25",X"4F",X"31",
		X"4F",X"3C",X"4F",X"47",X"4F",X"52",X"4F",X"77",X"4F",X"87",X"4F",X"B3",X"4F",X"CA",X"4F",X"E4",
		X"50",X"02",X"50",X"19",X"50",X"32",X"50",X"3C",X"50",X"68",X"50",X"82",X"50",X"89",X"50",X"9D",
		X"50",X"B7",X"50",X"DA",X"50",X"EB",X"51",X"02",X"51",X"23",X"51",X"31",X"51",X"42",X"4D",X"5C",
		X"4D",X"38",X"4D",X"4A",X"4C",X"EE",X"4C",X"99",X"4C",X"B5",X"4C",X"75",X"4C",X"88",X"4C",X"4C",
		X"4C",X"38",X"4C",X"2D",X"4C",X"10",X"4C",X"16",X"4C",X"20",X"4B",X"EC",X"1E",X"19",X"0A",X"10",
		X"13",X"11",X"12",X"1E",X"0A",X"1E",X"12",X"0F",X"0A",X"12",X"19",X"1E",X"0A",X"0B",X"18",X"0E",
		X"0A",X"1C",X"1F",X"1E",X"12",X"16",X"0F",X"1D",X"1D",X"0A",X"1D",X"19",X"1F",X"16",X"1D",X"AE",
		X"0A",X"1D",X"19",X"1F",X"16",X"9D",X"0F",X"16",X"13",X"17",X"13",X"18",X"0B",X"1E",X"0F",X"8E",
		X"1E",X"13",X"17",X"0F",X"1D",X"0A",X"03",X"2D",X"00",X"00",X"00",X"0A",X"A6",X"0D",X"19",X"0D",
		X"19",X"19",X"18",X"0A",X"21",X"0B",X"20",X"8F",X"0B",X"16",X"16",X"19",X"21",X"0A",X"02",X"0A",
		X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"0C",X"1F",X"23",X"13",X"98",X"0E",X"0F",X"1D",X"1E",
		X"1C",X"19",X"23",X"0A",X"1E",X"0B",X"18",X"15",X"19",X"20",X"1D",X"0A",X"1E",X"1C",X"0F",X"0B",
		X"0E",X"1D",X"0A",X"10",X"1C",X"19",X"17",X"0A",X"0B",X"0A",X"16",X"19",X"21",X"0F",X"1C",X"0A",
		X"16",X"0F",X"20",X"0F",X"96",X"0A",X"1D",X"19",X"1F",X"16",X"1D",X"0A",X"12",X"0B",X"20",X"0F",
		X"0A",X"0F",X"1D",X"0D",X"0B",X"1A",X"0F",X"8E",X"0A",X"1D",X"19",X"1F",X"16",X"0A",X"12",X"0B",
		X"1D",X"0A",X"0F",X"1D",X"0D",X"0B",X"1A",X"0F",X"8E",X"13",X"18",X"1D",X"0F",X"1C",X"1E",X"0A",
		X"0D",X"19",X"13",X"18",X"0A",X"1E",X"19",X"0A",X"0D",X"19",X"18",X"1E",X"13",X"18",X"1F",X"0F",
		X"0A",X"1A",X"16",X"0B",X"A3",X"1A",X"1C",X"0F",X"1D",X"1D",X"0A",X"1D",X"1E",X"0B",X"1C",X"1E",
		X"0A",X"1E",X"19",X"0A",X"0D",X"19",X"18",X"1E",X"13",X"18",X"1F",X"0F",X"0A",X"1A",X"16",X"0B",
		X"A3",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"0C",X"1F",X"23",X"27",X"13",X"98",X"0F",X"22",X"1E",
		X"1C",X"0B",X"0A",X"16",X"13",X"10",X"0F",X"0A",X"0F",X"20",X"0F",X"1C",X"23",X"8A",X"2D",X"00",
		X"00",X"80",X"0C",X"0F",X"21",X"0B",X"1C",X"0F",X"0A",X"19",X"10",X"0A",X"1E",X"12",X"0F",X"0A",
		X"12",X"13",X"11",X"12",X"0F",X"1C",X"0A",X"16",X"0F",X"20",X"0F",X"16",X"1D",X"AD",X"0B",X"18",
		X"23",X"19",X"18",X"0F",X"0A",X"0C",X"0F",X"16",X"19",X"21",X"0A",X"23",X"19",X"1F",X"0A",X"0D",
		X"0B",X"98",X"1E",X"0B",X"15",X"0F",X"0A",X"0B",X"0E",X"20",X"0B",X"18",X"1E",X"0B",X"11",X"0F",
		X"0A",X"19",X"10",X"0A",X"23",X"19",X"1F",X"AE",X"11",X"0B",X"17",X"0F",X"0A",X"19",X"20",X"0F",
		X"1C",X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"81",X"11",X"0B",X"17",X"0F",X"0A",X"19",
		X"20",X"0F",X"1C",X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"82",X"12",X"0F",X"1C",X"0A",
		X"1D",X"0F",X"22",X"23",X"0A",X"10",X"16",X"13",X"11",X"12",X"1E",X"0A",X"21",X"13",X"16",X"16",
		X"0A",X"1E",X"1C",X"0B",X"18",X"1B",X"1F",X"13",X"16",X"13",X"24",X"0F",X"0A",X"23",X"19",X"1F",
		X"1C",X"0A",X"0F",X"18",X"0F",X"17",X"13",X"0F",X"1D",X"AE",X"23",X"19",X"1F",X"0A",X"0B",X"1C",
		X"0F",X"0A",X"0B",X"0A",X"0C",X"19",X"1C",X"18",X"0A",X"12",X"0F",X"1C",X"19",X"AD",X"23",X"19",
		X"1F",X"0A",X"21",X"13",X"16",X"16",X"0A",X"10",X"13",X"11",X"12",X"1E",X"0A",X"1E",X"19",X"0A",
		X"1D",X"1F",X"1C",X"20",X"13",X"20",X"8F",X"1E",X"12",X"0F",X"0A",X"0F",X"20",X"13",X"16",X"0A",
		X"21",X"19",X"1C",X"16",X"0E",X"1D",X"0A",X"19",X"10",X"0A",X"1E",X"12",X"0F",X"0A",X"11",X"1C",
		X"0B",X"18",X"0E",X"0A",X"16",X"13",X"24",X"0B",X"1C",X"0E",X"AE",X"1E",X"19",X"0A",X"17",X"19",
		X"20",X"0F",X"0A",X"1F",X"1D",X"0F",X"0A",X"1E",X"12",X"0F",X"0A",X"1C",X"1F",X"18",X"0A",X"14",
		X"19",X"23",X"1D",X"1E",X"13",X"0D",X"15",X"AE",X"1E",X"0B",X"15",X"0F",X"0A",X"0D",X"0B",X"1C",
		X"0F",X"10",X"1F",X"16",X"16",X"0A",X"0B",X"13",X"17",X"AD",X"1E",X"12",X"0F",X"18",X"0A",X"10",
		X"13",X"1C",X"0F",X"0A",X"23",X"19",X"1F",X"1C",X"0A",X"16",X"0B",X"1D",X"0F",X"1C",X"0A",X"0B",
		X"1E",X"0A",X"0B",X"16",X"16",X"0A",X"0F",X"18",X"0F",X"17",X"13",X"0F",X"1D",X"AE",X"23",X"19",
		X"1F",X"0A",X"0D",X"0B",X"18",X"0A",X"19",X"18",X"16",X"23",X"0A",X"10",X"13",X"1C",X"0F",X"0A",
		X"13",X"18",X"0A",X"04",X"0A",X"0E",X"13",X"1C",X"0F",X"0D",X"1E",X"13",X"19",X"18",X"1D",X"AE",
		X"23",X"19",X"1F",X"0A",X"0E",X"19",X"0A",X"18",X"19",X"1E",X"0A",X"16",X"19",X"1D",X"0F",X"0A",
		X"0B",X"0A",X"16",X"13",X"10",X"0F",X"AD",X"13",X"10",X"0A",X"23",X"19",X"1F",X"1C",X"0A",X"1A",
		X"0B",X"1C",X"1E",X"18",X"0F",X"1C",X"0A",X"1D",X"12",X"19",X"19",X"1E",X"1D",X"0A",X"23",X"19",
		X"1F",X"AE",X"0C",X"1F",X"1E",X"0A",X"23",X"19",X"1F",X"0A",X"21",X"13",X"16",X"16",X"0A",X"16",
		X"19",X"1D",X"0F",X"0A",X"0B",X"0A",X"16",X"13",X"10",X"0F",X"AD",X"13",X"10",X"0A",X"23",X"19",
		X"1F",X"1C",X"0A",X"0F",X"18",X"0F",X"17",X"13",X"0F",X"1D",X"0A",X"1D",X"12",X"19",X"19",X"1E",
		X"0A",X"23",X"19",X"1F",X"AE",X"0B",X"10",X"1E",X"0F",X"1C",X"0A",X"23",X"19",X"1F",X"0A",X"0B",
		X"1C",X"0F",X"0A",X"0C",X"19",X"1C",X"18",X"AD",X"23",X"19",X"1F",X"0A",X"12",X"0B",X"20",X"0F",
		X"0A",X"1E",X"0F",X"17",X"1A",X"19",X"1C",X"0B",X"1C",X"23",X"0A",X"13",X"17",X"17",X"1F",X"18",
		X"13",X"1E",X"A3",X"1F",X"18",X"1E",X"13",X"16",X"0A",X"23",X"19",X"1F",X"0A",X"17",X"19",X"20",
		X"0F",X"0A",X"19",X"1C",X"0A",X"23",X"19",X"1F",X"1C",X"0A",X"0D",X"1C",X"0F",X"0B",X"1E",X"13",
		X"19",X"18",X"0A",X"13",X"1D",X"0A",X"0D",X"19",X"17",X"1A",X"16",X"0F",X"1E",X"0F",X"AE",X"12",
		X"0F",X"1C",X"0F",X"0A",X"0B",X"1C",X"0F",X"0A",X"23",X"19",X"1F",X"1C",X"0A",X"0F",X"18",X"0F",
		X"17",X"13",X"0F",X"1D",X"AE",X"1E",X"12",X"0F",X"0A",X"0D",X"23",X"0D",X"16",X"19",X"1A",X"1D",
		X"B2",X"0E",X"19",X"12",X"1C",X"1E",X"0A",X"2A",X"05",X"00",X"00",X"AB",X"24",X"19",X"12",X"1C",
		X"1E",X"0A",X"2A",X"07",X"00",X"00",X"AB",X"17",X"19",X"12",X"1C",X"1E",X"0A",X"2A",X"09",X"00",
		X"00",X"AB",X"0B",X"10",X"1E",X"0F",X"1C",X"0A",X"23",X"19",X"1F",X"0A",X"1D",X"12",X"19",X"19",
		X"1E",X"0A",X"1E",X"12",X"0F",X"17",X"0A",X"21",X"13",X"1E",X"12",X"0A",X"23",X"19",X"1F",X"1C",
		X"0A",X"16",X"0B",X"1D",X"0F",X"1C",X"AD",X"1E",X"0B",X"11",X"0A",X"1E",X"12",X"0F",X"13",X"1C",
		X"0A",X"1D",X"19",X"1F",X"16",X"1D",X"AD",X"19",X"1C",X"0A",X"10",X"19",X"16",X"16",X"19",X"21",
		X"0A",X"1E",X"12",X"0F",X"17",X"0A",X"13",X"18",X"1E",X"19",X"0A",X"1E",X"12",X"0F",X"0A",X"11",
		X"1C",X"0B",X"18",X"0E",X"0A",X"16",X"13",X"24",X"0B",X"1C",X"0E",X"2C",X"1D",X"0A",X"17",X"19",
		X"1F",X"1E",X"92",X"10",X"19",X"1C",X"0A",X"0F",X"22",X"1E",X"1C",X"0B",X"0A",X"0C",X"19",X"18",
		X"1F",X"1D",X"0A",X"1A",X"19",X"13",X"18",X"1E",X"1D",X"AE",X"0E",X"19",X"0A",X"18",X"19",X"1E",
		X"0A",X"16",X"0F",X"1E",X"0A",X"01",X"03",X"0A",X"1D",X"19",X"1F",X"16",X"1D",X"0A",X"0F",X"1D",
		X"0D",X"0B",X"1A",X"8F",X"13",X"18",X"1E",X"19",X"0A",X"1E",X"12",X"0F",X"0A",X"11",X"1C",X"0B",
		X"18",X"0E",X"0A",X"16",X"13",X"24",X"0B",X"1C",X"0E",X"2C",X"1D",X"0A",X"17",X"19",X"1F",X"1E",
		X"12",X"AD",X"10",X"19",X"1C",X"0A",X"1E",X"12",X"0F",X"23",X"0A",X"21",X"13",X"16",X"16",X"0A",
		X"12",X"0B",X"1F",X"18",X"1E",X"0A",X"23",X"19",X"9F",X"13",X"18",X"0A",X"1E",X"12",X"0F",X"13",
		X"1C",X"0A",X"1C",X"0F",X"0E",X"0A",X"12",X"19",X"1E",X"0A",X"13",X"18",X"10",X"0F",X"1C",X"18",
		X"19",X"AE",X"1E",X"12",X"0F",X"0A",X"18",X"23",X"17",X"1A",X"12",X"B2",X"21",X"13",X"1E",X"12",
		X"0A",X"0B",X"0A",X"0D",X"0B",X"1A",X"1E",X"1F",X"1C",X"0F",X"0E",X"0A",X"1D",X"19",X"1F",X"16",
		X"2D",X"0A",X"23",X"19",X"1F",X"0A",X"11",X"13",X"20",X"0F",X"0A",X"16",X"13",X"10",X"0F",X"0A",
		X"0B",X"18",X"0E",X"0A",X"10",X"1C",X"0F",X"8F",X"1E",X"12",X"0F",X"0A",X"18",X"23",X"17",X"1A",
		X"12",X"0A",X"16",X"19",X"0D",X"15",X"0F",X"0E",X"0A",X"13",X"18",X"0A",X"1D",X"1E",X"19",X"18",
		X"0F",X"AE",X"1E",X"0B",X"18",X"15",X"19",X"20",X"B2",X"23",X"19",X"1F",X"0A",X"17",X"1F",X"1D",
		X"1E",X"0A",X"0E",X"0F",X"1D",X"1E",X"1C",X"19",X"23",X"0A",X"12",X"13",X"9D",X"1E",X"1C",X"0F",
		X"0B",X"0E",X"1D",X"0A",X"10",X"1C",X"19",X"17",X"0A",X"0B",X"0A",X"16",X"19",X"21",X"0F",X"1C",
		X"0A",X"16",X"0F",X"20",X"0F",X"16",X"AD",X"0B",X"18",X"0E",X"0A",X"12",X"13",X"1D",X"0A",X"1E",
		X"1F",X"1C",X"1C",X"0F",X"1E",X"0A",X"10",X"1C",X"19",X"17",X"0A",X"1E",X"12",X"0F",X"0A",X"1D",
		X"0B",X"17",X"0F",X"0A",X"16",X"0F",X"20",X"0F",X"16",X"AE",X"13",X"10",X"0A",X"23",X"19",X"1F",
		X"0A",X"17",X"1F",X"1D",X"1E",X"0A",X"1A",X"0B",X"18",X"13",X"8D",X"1D",X"1E",X"0F",X"1A",X"0A",
		X"19",X"18",X"0A",X"1E",X"12",X"0F",X"0A",X"16",X"0B",X"1F",X"18",X"0D",X"12",X"0A",X"1A",X"0B",
		X"0E",X"AD",X"13",X"1E",X"0A",X"21",X"13",X"16",X"16",X"0A",X"0F",X"14",X"0F",X"0D",X"1E",X"0A",
		X"23",X"19",X"1F",X"0A",X"19",X"1F",X"1E",X"0A",X"19",X"10",X"0A",X"1E",X"1C",X"19",X"1F",X"0C",
		X"16",X"0F",X"AE",X"1E",X"12",X"0F",X"0A",X"0C",X"19",X"19",X"17",X"0A",X"0C",X"13",X"1C",X"0E",
		X"B2",X"12",X"0F",X"0A",X"1A",X"0B",X"1E",X"1C",X"19",X"16",X"1D",X"0A",X"0B",X"0C",X"19",X"20",
		X"0F",X"AD",X"0B",X"18",X"0E",X"0A",X"19",X"18",X"16",X"23",X"0A",X"0B",X"0A",X"10",X"0F",X"21",
		X"0A",X"15",X"18",X"19",X"21",X"0A",X"12",X"19",X"21",X"0A",X"1E",X"19",X"0A",X"0E",X"0F",X"0B",
		X"16",X"0A",X"21",X"13",X"1E",X"12",X"0A",X"12",X"13",X"17",X"AE",X"0E",X"19",X"12",X"1C",X"1E",
		X"0A",X"21",X"0B",X"20",X"8F",X"24",X"19",X"12",X"1C",X"1E",X"0A",X"21",X"0B",X"20",X"8F",X"17",
		X"19",X"12",X"1C",X"1E",X"0A",X"21",X"0B",X"20",X"8F",X"21",X"0B",X"20",X"0F",X"0A",X"1A",X"19",
		X"13",X"18",X"1E",X"9D",X"0C",X"19",X"18",X"1F",X"1D",X"0A",X"1A",X"0F",X"1C",X"0D",X"0F",X"18",
		X"9E",X"0C",X"19",X"18",X"1F",X"1D",X"0A",X"1A",X"19",X"13",X"18",X"1E",X"9D",X"1A",X"1C",X"0F",
		X"1D",X"1D",X"8A",X"31",X"1D",X"13",X"18",X"11",X"16",X"0F",X"0A",X"1A",X"16",X"0B",X"23",X"B1",
		X"0A",X"1E",X"19",X"0A",X"1D",X"1E",X"0B",X"1C",X"9E",X"19",X"9C",X"13",X"18",X"1D",X"0F",X"1C",
		X"1E",X"0A",X"0B",X"0E",X"0E",X"13",X"1E",X"13",X"19",X"18",X"0B",X"16",X"0A",X"0D",X"19",X"13",
		X"18",X"1D",X"0A",X"10",X"19",X"9C",X"1C",X"0F",X"0B",X"0E",X"23",X"0A",X"10",X"19",X"1C",X"8A",
		X"31",X"0E",X"1F",X"0B",X"16",X"0A",X"1A",X"16",X"0B",X"23",X"B1",X"0C",X"19",X"19",X"17",X"0A",
		X"0C",X"13",X"1C",X"0E",X"0A",X"21",X"0B",X"20",X"8F",X"1E",X"0B",X"18",X"15",X"19",X"20",X"0A",
		X"21",X"0B",X"20",X"8F",X"13",X"18",X"10",X"0F",X"1C",X"18",X"19",X"0A",X"21",X"0B",X"20",X"8F",
		X"1A",X"1C",X"0F",X"1A",X"0B",X"1C",X"0F",X"0A",X"1E",X"19",X"0A",X"0E",X"0F",X"10",X"0F",X"18",
		X"0E",X"0A",X"1E",X"12",X"23",X"0A",X"1D",X"0F",X"16",X"90",X"0D",X"1F",X"1D",X"1E",X"19",X"97",
		X"13",X"18",X"10",X"0F",X"1C",X"18",X"99",X"1E",X"12",X"23",X"0A",X"11",X"0B",X"17",X"0F",X"0A",
		X"13",X"1D",X"0A",X"19",X"20",X"0F",X"9C",X"13",X"18",X"13",X"1E",X"13",X"0B",X"16",X"0A",X"1E",
		X"0F",X"1D",X"1E",X"1D",X"0A",X"13",X"18",X"0E",X"13",X"0D",X"0B",X"1E",X"8F",X"0B",X"16",X"16",
		X"0A",X"1D",X"23",X"1D",X"1E",X"0F",X"17",X"1D",X"0A",X"11",X"99",X"1C",X"0B",X"17",X"0A",X"0F",
		X"1C",X"1C",X"19",X"1C",X"8A",X"1C",X"19",X"17",X"0A",X"0F",X"1C",X"1C",X"19",X"1C",X"8A",X"1C",
		X"0B",X"17",X"0A",X"1E",X"0F",X"1D",X"1E",X"0A",X"10",X"19",X"16",X"16",X"19",X"21",X"9D",X"1A",
		X"1C",X"0F",X"1D",X"1D",X"0A",X"0B",X"0E",X"20",X"0B",X"18",X"0D",X"0F",X"0A",X"1E",X"19",X"0A",
		X"0F",X"22",X"13",X"9E",X"1C",X"0B",X"17",X"0A",X"0F",X"1C",X"1C",X"19",X"1C",X"1D",X"0A",X"0E",
		X"0F",X"1E",X"0F",X"0D",X"1E",X"0F",X"8E",X"18",X"19",X"8A",X"18",X"19",X"0A",X"0D",X"17",X"19",
		X"1D",X"8A",X"0D",X"17",X"19",X"1D",X"0A",X"1C",X"0B",X"17",X"0A",X"0F",X"1C",X"1C",X"19",X"9C",
		X"10",X"1C",X"19",X"18",X"1E",X"0A",X"0E",X"19",X"19",X"1C",X"0A",X"17",X"1F",X"1D",X"1E",X"0A",
		X"0C",X"0F",X"0A",X"19",X"1A",X"0F",X"98",X"19",X"1C",X"0A",X"1E",X"0B",X"0C",X"16",X"0F",X"0A",
		X"1E",X"19",X"1A",X"0A",X"1C",X"0B",X"1D",X"13",X"0F",X"0E",X"0A",X"10",X"19",X"1C",X"0A",X"1E",
		X"0F",X"1D",X"9E",X"19",X"1C",X"0A",X"21",X"1C",X"13",X"1E",X"0F",X"0A",X"1A",X"1C",X"19",X"1E",
		X"0F",X"0D",X"1E",X"0A",X"10",X"0B",X"13",X"16",X"1F",X"1C",X"8F",X"1D",X"21",X"13",X"1E",X"0D",
		X"12",X"0A",X"1E",X"0F",X"1D",X"9E",X"0B",X"1F",X"1E",X"19",X"0A",X"1F",X"9A",X"0B",X"0E",X"20",
		X"0B",X"18",X"0D",X"8F",X"1C",X"13",X"11",X"12",X"1E",X"0A",X"0D",X"19",X"13",X"98",X"12",X"13",
		X"11",X"12",X"0A",X"1D",X"0D",X"19",X"1C",X"0F",X"0A",X"1C",X"0F",X"1D",X"0F",X"9E",X"16",X"0F",
		X"10",X"1E",X"0A",X"0D",X"19",X"13",X"98",X"0D",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"0D",X"19",
		X"13",X"98",X"1D",X"16",X"0B",X"17",X"0A",X"1D",X"21",X"13",X"1E",X"0D",X"92",X"19",X"18",X"0F",
		X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"1D",X"1E",X"0B",X"1C",X"9E",X"1E",X"21",X"19",
		X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"1D",X"1E",X"0B",X"1C",X"9E",X"1D",X"19",X"1F",
		X"18",X"0E",X"0A",X"16",X"13",X"18",X"8F",X"0C",X"19",X"19",X"15",X"15",X"0F",X"0F",X"1A",X"13",
		X"18",X"11",X"0A",X"1E",X"19",X"1E",X"0B",X"16",X"1D",X"8A",X"16",X"0F",X"10",X"1E",X"0A",X"1D",
		X"16",X"19",X"1E",X"0A",X"0D",X"19",X"13",X"18",X"9D",X"0D",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",
		X"1D",X"16",X"19",X"1E",X"0A",X"0D",X"19",X"13",X"18",X"9D",X"1C",X"13",X"11",X"12",X"1E",X"0A",
		X"1D",X"16",X"19",X"1E",X"0A",X"0D",X"19",X"13",X"18",X"9D",X"1A",X"0B",X"13",X"0E",X"0A",X"0D",
		X"1C",X"0F",X"0E",X"13",X"1E",X"9D",X"10",X"1C",X"0F",X"0F",X"0A",X"17",X"0F",X"98",X"1E",X"19",
		X"1E",X"0B",X"16",X"0A",X"1E",X"13",X"17",X"0F",X"0A",X"13",X"18",X"0A",X"17",X"13",X"18",X"1F",
		X"1E",X"0F",X"9D",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"17",X"0F",X"18",X"0A",X"1A",X"16",X"0B",
		X"23",X"0F",X"8E",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"1D",X"13",X"18",X"11",X"16",X"0F",X"0A",
		X"1A",X"16",X"0B",X"23",X"0F",X"9C",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"0E",X"1F",X"0B",X"16",
		X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"9C",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"0D",X"1C",X"0F",
		X"0E",X"13",X"1E",X"1D",X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"8E",X"0B",X"20",X"0F",X"1C",X"0B",
		X"11",X"0F",X"0A",X"1E",X"13",X"17",X"0F",X"0A",X"1A",X"0F",X"1C",X"0A",X"0D",X"1C",X"0F",X"0E",
		X"13",X"9E",X"11",X"0B",X"17",X"0F",X"0A",X"0B",X"0E",X"14",X"1F",X"1D",X"1E",X"17",X"0F",X"18",
		X"1E",X"1D",X"8A",X"17",X"0F",X"18",X"0A",X"10",X"19",X"1C",X"0A",X"01",X"0A",X"0D",X"1C",X"0F",
		X"0E",X"13",X"1E",X"0A",X"11",X"0B",X"17",X"8F",X"12",X"13",X"11",X"12",X"0A",X"1D",X"0D",X"19",
		X"1C",X"0F",X"0A",X"1E",X"19",X"0A",X"0E",X"0B",X"1E",X"0F",X"0A",X"0B",X"16",X"16",X"19",X"21",
		X"0F",X"8E",X"1A",X"1C",X"13",X"0D",X"13",X"18",X"11",X"0A",X"1D",X"0F",X"16",X"0F",X"0D",X"1E",
		X"13",X"19",X"98",X"16",X"0F",X"10",X"1E",X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"1F",X"18",X"13",
		X"1E",X"9D",X"0D",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"1F",X"18",
		X"13",X"1E",X"9D",X"1C",X"13",X"11",X"12",X"1E",X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"1F",X"18",
		X"13",X"1E",X"9D",X"1F",X"18",X"13",X"1E",X"1D",X"0A",X"1C",X"0F",X"1B",X"1F",X"13",X"1C",X"0F",
		X"0E",X"0A",X"10",X"19",X"1C",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"1F",X"18",X"13",X"1E",
		X"1D",X"0A",X"1C",X"0F",X"1B",X"1F",X"13",X"1C",X"0F",X"0E",X"0A",X"10",X"19",X"1C",X"0A",X"0C",
		X"19",X"18",X"1F",X"1D",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"17",X"13",X"18",X"13",X"17",
		X"1F",X"17",X"0A",X"1F",X"18",X"13",X"1E",X"1D",X"0A",X"10",X"19",X"1C",X"0A",X"0B",X"18",X"23",
		X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"0E",X"13",X"10",X"10",X"13",X"0D",X"1F",X"16",X"1E",
		X"23",X"0A",X"19",X"10",X"0A",X"1A",X"16",X"0B",X"A3",X"16",X"0F",X"1E",X"1E",X"0F",X"1C",X"1D",
		X"0A",X"10",X"19",X"1C",X"0A",X"12",X"13",X"11",X"12",X"0F",X"1D",X"1E",X"0A",X"1D",X"0D",X"19",
		X"1C",X"8F",X"1C",X"0F",X"1D",X"1E",X"19",X"1C",X"0F",X"0A",X"10",X"0B",X"0D",X"1E",X"19",X"1C",
		X"23",X"0A",X"1D",X"0F",X"1E",X"1E",X"13",X"18",X"11",X"9D",X"0D",X"16",X"0F",X"0B",X"1C",X"0A",
		X"0C",X"19",X"19",X"15",X"15",X"0F",X"0F",X"1A",X"13",X"18",X"11",X"0A",X"1E",X"19",X"1E",X"0B",
		X"16",X"9D",X"12",X"13",X"11",X"12",X"0A",X"1D",X"0D",X"19",X"1C",X"0F",X"0A",X"1E",X"0B",X"0C",
		X"16",X"0F",X"0A",X"1C",X"0F",X"1D",X"0F",X"9E",X"0B",X"1F",X"1E",X"19",X"0A",X"0D",X"23",X"0D",
		X"16",X"8F",X"1D",X"0F",X"1E",X"0A",X"0B",X"1E",X"1E",X"1C",X"0B",X"0D",X"1E",X"0A",X"17",X"19",
		X"0E",X"0F",X"0A",X"17",X"0F",X"1D",X"1D",X"0B",X"11",X"8F",X"1D",X"0F",X"1E",X"0A",X"12",X"13",
		X"11",X"12",X"0F",X"1D",X"1E",X"0A",X"1D",X"0D",X"19",X"1C",X"0F",X"0A",X"18",X"0B",X"17",X"8F",
		X"1F",X"1D",X"0F",X"0A",X"2C",X"1C",X"1F",X"18",X"2C",X"0A",X"1E",X"19",X"0A",X"1D",X"0F",X"16",
		X"0F",X"0D",X"1E",X"8A",X"1F",X"1D",X"0F",X"0A",X"2C",X"0B",X"13",X"17",X"2C",X"0A",X"1E",X"19",
		X"0A",X"0D",X"12",X"0B",X"18",X"11",X"0F",X"0A",X"1E",X"12",X"0F",X"0A",X"20",X"0B",X"16",X"1F",
		X"8F",X"23",X"0F",X"9D",X"0B",X"0E",X"14",X"1F",X"1D",X"1E",X"17",X"0F",X"18",X"9E",X"16",X"0F",
		X"1E",X"1E",X"0F",X"9C",X"1F",X"1D",X"0F",X"0A",X"2C",X"0B",X"13",X"17",X"2C",X"0A",X"1E",X"19",
		X"0A",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"16",X"0F",X"1E",X"1E",X"0F",X"9C",X"0A",X"10",X"0B",
		X"13",X"16",X"1F",X"1C",X"8F",X"10",X"0B",X"0D",X"1E",X"19",X"1C",X"23",X"0A",X"1D",X"0F",X"1E",
		X"1E",X"13",X"18",X"11",X"1D",X"0A",X"1C",X"0F",X"1D",X"1E",X"19",X"1C",X"0F",X"8E",X"0C",X"23",
		X"0A",X"19",X"1A",X"0F",X"18",X"13",X"18",X"11",X"0A",X"10",X"1C",X"19",X"18",X"1E",X"0A",X"0E",
		X"19",X"19",X"1C",X"0A",X"19",X"1C",X"0A",X"1E",X"0B",X"0C",X"16",X"0F",X"0A",X"1E",X"19",X"9A",
		X"0B",X"18",X"0E",X"0A",X"1E",X"1F",X"1C",X"18",X"13",X"18",X"11",X"0A",X"11",X"0B",X"17",X"0F",
		X"0A",X"19",X"18",X"0A",X"0B",X"18",X"0E",X"0A",X"19",X"10",X"90",X"0A",X"0D",X"16",X"0F",X"0B",
		X"1C",X"0F",X"8E",X"12",X"13",X"11",X"12",X"0A",X"1D",X"0D",X"19",X"1C",X"0F",X"0A",X"1E",X"0B",
		X"0C",X"16",X"0F",X"0A",X"1C",X"0F",X"1D",X"0F",X"9E",X"0E",X"0B",X"13",X"16",X"23",X"0A",X"17",
		X"0B",X"1C",X"15",X"1D",X"17",X"0B",X"98",X"0F",X"1E",X"0F",X"1C",X"18",X"0B",X"16",X"0A",X"12",
		X"0F",X"1C",X"19",X"2C",X"9D",X"0D",X"1C",X"0F",X"0E",X"13",X"1E",X"1D",X"8A",X"1F",X"1D",X"0F",
		X"0A",X"2C",X"0B",X"13",X"17",X"2C",X"0A",X"1E",X"19",X"0A",X"0D",X"0F",X"18",X"1E",X"0F",X"9C",
		X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"16",X"13",X"18",X"0F",X"0A",X"0C",X"23",X"0A",X"1A",X"1C",
		X"0F",X"1D",X"1D",X"13",X"18",X"11",X"0A",X"0B",X"0E",X"20",X"0B",X"18",X"0D",X"8F",X"0F",X"18",
		X"1E",X"0F",X"1C",X"0A",X"1E",X"12",X"23",X"0A",X"18",X"0B",X"17",X"0F",X"0A",X"17",X"23",X"0A",
		X"16",X"19",X"1C",X"0E",X"A9",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"23",X"19",X"1F",X"1C",X"0A",
		X"13",X"18",X"13",X"1E",X"13",X"0B",X"16",X"9D",X"11",X"19",X"19",X"0E",X"0A",X"1D",X"12",X"19",
		X"19",X"1E",X"13",X"18",X"91",X"17",X"0B",X"22",X"13",X"17",X"1F",X"17",X"0A",X"05",X"0A",X"0F",
		X"18",X"1E",X"1C",X"23",X"9D",X"1F",X"1D",X"0F",X"0A",X"27",X"1C",X"1F",X"18",X"27",X"0A",X"1E",
		X"19",X"0A",X"1D",X"0F",X"16",X"0F",X"0D",X"1E",X"0A",X"16",X"0F",X"1E",X"1E",X"0F",X"1C",X"0A",
		X"0A",X"0A",X"0A",X"27",X"0B",X"13",X"17",X"27",X"0A",X"1E",X"19",X"0A",X"0F",X"18",X"1E",X"0F",
		X"1C",X"0A",X"16",X"0F",X"1E",X"1E",X"0F",X"9C",X"2A",X"0D",X"2B",X"0A",X"01",X"09",X"08",X"04",
		X"0A",X"21",X"13",X"16",X"16",X"13",X"0B",X"17",X"1D",X"0A",X"0F",X"16",X"0F",X"0D",X"1E",X"1C",
		X"19",X"18",X"13",X"0D",X"1D",X"0A",X"13",X"18",X"0D",X"AE",X"11",X"0B",X"17",X"0F",X"0A",X"19",
		X"20",X"0F",X"9C",X"10",X"1C",X"0F",X"0F",X"0A",X"1A",X"16",X"0B",X"A3",X"1E",X"12",X"13",X"1D",
		X"0A",X"13",X"1D",X"0A",X"13",X"18",X"10",X"0F",X"1C",X"18",X"99",X"0E",X"0F",X"1D",X"13",X"11",
		X"18",X"0F",X"0E",X"0A",X"0C",X"23",X"0A",X"21",X"13",X"16",X"16",X"13",X"0B",X"17",X"1D",X"0A",
		X"0F",X"16",X"0F",X"0D",X"1E",X"1C",X"19",X"18",X"13",X"0D",X"1D",X"0A",X"13",X"18",X"0D",X"AE",
		X"0B",X"16",X"16",X"0A",X"1C",X"13",X"11",X"12",X"1E",X"1D",X"0A",X"1C",X"0F",X"1D",X"0F",X"1C",
		X"20",X"0F",X"8E",X"1C",X"1F",X"18",X"0A",X"1F",X"1A",X"27",X"1C",X"13",X"11",X"12",X"9E",X"1C",
		X"1F",X"18",X"0A",X"1F",X"1A",X"27",X"16",X"0F",X"10",X"9E",X"1C",X"1F",X"18",X"0A",X"0E",X"19",
		X"21",X"18",X"27",X"1C",X"13",X"11",X"12",X"9E",X"1C",X"1F",X"18",X"0A",X"0E",X"19",X"21",X"18",
		X"27",X"16",X"0F",X"10",X"9E",X"0B",X"13",X"17",X"0A",X"1F",X"1A",X"27",X"1C",X"13",X"11",X"12",
		X"9E",X"0B",X"13",X"17",X"0A",X"1F",X"1A",X"27",X"16",X"0F",X"10",X"9E",X"0B",X"13",X"17",X"0A",
		X"0E",X"19",X"21",X"18",X"27",X"1C",X"13",X"11",X"12",X"9E",X"0B",X"13",X"17",X"0A",X"0E",X"19",
		X"21",X"18",X"27",X"16",X"0F",X"10",X"9E",X"1E",X"1C",X"13",X"11",X"11",X"0F",X"9C",X"58",X"A4",
		X"58",X"AC",X"58",X"B4",X"58",X"BC",X"58",X"C0",X"58",X"D0",X"58",X"D4",X"58",X"D8",X"58",X"DC",
		X"58",X"EC",X"58",X"FC",X"59",X"10",X"59",X"14",X"59",X"1C",X"59",X"20",X"59",X"28",X"59",X"38",
		X"59",X"48",X"59",X"60",X"36",X"CC",X"05",X"11",X"2E",X"DC",X"86",X"11",X"2A",X"80",X"08",X"99",
		X"00",X"00",X"87",X"99",X"21",X"80",X"09",X"99",X"00",X"00",X"87",X"99",X"36",X"80",X"8A",X"22",
		X"36",X"80",X"0A",X"22",X"28",X"90",X"0D",X"22",X"17",X"A0",X"0B",X"99",X"17",X"A8",X"8C",X"99",
		X"3A",X"20",X"8E",X"88",X"2F",X"10",X"9F",X"99",X"2F",X"10",X"AC",X"99",X"23",X"D7",X"3F",X"BB",
		X"00",X"00",X"42",X"BB",X"25",X"DF",X"40",X"44",X"34",X"E7",X"86",X"11",X"28",X"16",X"3D",X"BB",
		X"16",X"C0",X"3F",X"33",X"00",X"00",X"43",X"33",X"20",X"D0",X"C4",X"33",X"30",X"80",X"42",X"22",
		X"00",X"00",X"45",X"22",X"27",X"A0",X"39",X"22",X"19",X"B0",X"47",X"22",X"23",X"C0",X"C8",X"22",
		X"21",X"80",X"C6",X"99",X"24",X"60",X"1F",X"33",X"00",X"00",X"C9",X"33",X"2A",X"40",X"CA",X"88",
		X"3A",X"2A",X"4B",X"11",X"31",X"60",X"CC",X"22",X"28",X"16",X"3E",X"BB",X"16",X"C0",X"3F",X"33",
		X"00",X"00",X"43",X"33",X"20",X"D0",X"C4",X"33",X"10",X"30",X"50",X"11",X"10",X"40",X"51",X"11",
		X"10",X"50",X"58",X"11",X"10",X"60",X"D2",X"11",X"24",X"57",X"65",X"11",X"00",X"00",X"66",X"55",
		X"00",X"00",X"67",X"11",X"49",X"77",X"68",X"11",X"26",X"97",X"69",X"11",X"3D",X"A7",X"EB",X"77",
		X"2E",X"77",X"6A",X"11",X"00",X"00",X"EB",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"34",X"40",X"33",X"48",X"C6",X"11",X"BD",X"E0",X"72",X"84",X"0F",X"4C",X"A7",X"44",X"33",X"45",
		X"5A",X"26",X"F3",X"35",X"C0",X"33",X"48",X"C6",X"11",X"34",X"04",X"8D",X"09",X"33",X"45",X"6A",
		X"E4",X"26",X"F8",X"35",X"84",X"39",X"E6",X"44",X"27",X"4A",X"6A",X"44",X"26",X"F7",X"BD",X"E0",
		X"72",X"49",X"C6",X"70",X"3D",X"8B",X"0C",X"84",X"FE",X"C6",X"93",X"1F",X"01",X"30",X"89",X"FE",
		X"00",X"30",X"89",X"02",X"00",X"8C",X"7C",X"00",X"25",X"04",X"30",X"89",X"90",X"00",X"86",X"00",
		X"BD",X"E0",X"83",X"85",X"F0",X"27",X"EA",X"85",X"0F",X"27",X"E6",X"5D",X"26",X"E3",X"1F",X"10",
		X"A7",X"C4",X"BD",X"E0",X"72",X"84",X"07",X"8B",X"02",X"A7",X"42",X"A7",X"43",X"86",X"8E",X"A7",
		X"41",X"7E",X"60",X"98",X"E6",X"41",X"C1",X"94",X"24",X"0D",X"6A",X"43",X"26",X"19",X"A6",X"42",
		X"A7",X"43",X"6C",X"41",X"7E",X"60",X"98",X"6C",X"41",X"E6",X"41",X"C1",X"BA",X"23",X"09",X"BD",
		X"E0",X"72",X"84",X"0F",X"4C",X"A7",X"44",X"39",X"34",X"01",X"1A",X"F0",X"10",X"8E",X"60",X"D4",
		X"8E",X"02",X"08",X"A6",X"C4",X"E6",X"41",X"C1",X"94",X"24",X"0A",X"C0",X"94",X"30",X"85",X"50",
		X"58",X"31",X"A5",X"C6",X"94",X"FD",X"C8",X"84",X"BF",X"C8",X"86",X"10",X"BF",X"C8",X"82",X"CB",
		X"08",X"C0",X"B9",X"23",X"08",X"50",X"CB",X"08",X"2B",X"08",X"F7",X"C8",X"87",X"86",X"02",X"B7",
		X"C8",X"80",X"35",X"81",X"00",X"00",X"02",X"00",X"02",X"00",X"32",X"30",X"32",X"30",X"22",X"20",
		X"22",X"20",X"02",X"00",X"30",X"4E",X"10",X"8E",X"61",X"05",X"CC",X"06",X"00",X"10",X"AF",X"02",
		X"E7",X"84",X"5C",X"6F",X"01",X"30",X"04",X"4A",X"26",X"F3",X"CC",X"62",X"FF",X"ED",X"1E",X"6F",
		X"48",X"CC",X"63",X"95",X"ED",X"4C",X"39",X"61",X"21",X"61",X"49",X"61",X"71",X"61",X"99",X"61",
		X"C1",X"61",X"E9",X"62",X"11",X"62",X"39",X"62",X"61",X"62",X"89",X"62",X"B1",X"62",X"D9",X"00",
		X"00",X"72",X"71",X"75",X"43",X"43",X"43",X"43",X"43",X"72",X"71",X"75",X"43",X"43",X"43",X"43",
		X"43",X"72",X"71",X"75",X"43",X"43",X"43",X"43",X"43",X"72",X"71",X"75",X"43",X"43",X"43",X"43",
		X"43",X"72",X"71",X"75",X"43",X"43",X"43",X"43",X"43",X"4E",X"53",X"75",X"43",X"43",X"43",X"43",
		X"43",X"4F",X"54",X"75",X"43",X"43",X"43",X"43",X"43",X"50",X"55",X"75",X"43",X"43",X"43",X"43",
		X"43",X"51",X"56",X"75",X"43",X"43",X"43",X"43",X"43",X"52",X"57",X"75",X"43",X"43",X"43",X"43",
		X"43",X"4E",X"58",X"76",X"75",X"43",X"43",X"43",X"43",X"4F",X"59",X"76",X"75",X"43",X"43",X"43",
		X"43",X"50",X"5A",X"76",X"75",X"43",X"43",X"43",X"43",X"51",X"5B",X"76",X"75",X"43",X"43",X"43",
		X"43",X"52",X"5C",X"76",X"75",X"43",X"43",X"43",X"43",X"4E",X"5D",X"62",X"75",X"43",X"43",X"43",
		X"43",X"4F",X"5E",X"63",X"75",X"43",X"43",X"43",X"43",X"50",X"5F",X"64",X"75",X"43",X"43",X"43",
		X"43",X"51",X"60",X"65",X"75",X"43",X"43",X"43",X"43",X"52",X"61",X"66",X"75",X"43",X"43",X"43",
		X"43",X"4E",X"5D",X"67",X"76",X"75",X"43",X"43",X"43",X"4F",X"5E",X"68",X"76",X"75",X"43",X"43",
		X"43",X"50",X"5F",X"69",X"76",X"75",X"43",X"43",X"43",X"51",X"60",X"6A",X"76",X"75",X"43",X"43",
		X"43",X"52",X"61",X"6B",X"76",X"75",X"43",X"43",X"43",X"4E",X"5D",X"6C",X"62",X"75",X"43",X"43",
		X"43",X"4F",X"5E",X"6D",X"63",X"75",X"43",X"43",X"43",X"50",X"5F",X"6E",X"64",X"75",X"43",X"43",
		X"43",X"51",X"60",X"6F",X"65",X"75",X"43",X"43",X"43",X"52",X"61",X"70",X"66",X"75",X"43",X"43",
		X"43",X"4E",X"5D",X"6C",X"67",X"76",X"75",X"43",X"43",X"4F",X"5E",X"6D",X"68",X"76",X"75",X"43",
		X"43",X"50",X"5F",X"6E",X"69",X"76",X"75",X"43",X"43",X"51",X"60",X"6F",X"6A",X"76",X"75",X"43",
		X"43",X"52",X"61",X"70",X"6B",X"76",X"75",X"43",X"43",X"4E",X"5D",X"6C",X"6C",X"62",X"75",X"43",
		X"43",X"4F",X"5E",X"6D",X"6D",X"63",X"75",X"43",X"43",X"50",X"5F",X"6E",X"6E",X"64",X"75",X"43",
		X"43",X"51",X"60",X"6F",X"6F",X"65",X"75",X"43",X"43",X"52",X"61",X"70",X"70",X"66",X"75",X"43",
		X"43",X"4E",X"5D",X"6C",X"6C",X"67",X"76",X"75",X"43",X"4F",X"5E",X"6D",X"6D",X"68",X"76",X"75",
		X"43",X"50",X"5F",X"6E",X"6E",X"69",X"76",X"75",X"43",X"51",X"60",X"6F",X"6F",X"6A",X"76",X"75",
		X"43",X"52",X"61",X"70",X"70",X"6B",X"76",X"75",X"43",X"4E",X"5D",X"6C",X"6C",X"6C",X"62",X"75",
		X"43",X"4F",X"5E",X"6D",X"6D",X"6D",X"63",X"75",X"43",X"50",X"5F",X"6E",X"6E",X"6E",X"64",X"75",
		X"43",X"51",X"60",X"6F",X"6F",X"6F",X"65",X"75",X"43",X"52",X"61",X"70",X"70",X"70",X"66",X"75",
		X"43",X"4E",X"5D",X"6C",X"6C",X"6C",X"67",X"76",X"75",X"4F",X"5E",X"6D",X"6D",X"6D",X"68",X"76",
		X"75",X"50",X"5F",X"6E",X"6E",X"6E",X"69",X"76",X"75",X"51",X"60",X"6F",X"6F",X"6F",X"6A",X"76",
		X"75",X"52",X"61",X"70",X"70",X"70",X"6B",X"76",X"75",X"4E",X"5D",X"6C",X"6C",X"6C",X"6C",X"62",
		X"75",X"4F",X"5E",X"6D",X"6D",X"6D",X"6D",X"63",X"75",X"50",X"5F",X"6E",X"6E",X"6E",X"6E",X"64",
		X"75",X"51",X"60",X"6F",X"6F",X"6F",X"6F",X"65",X"75",X"52",X"61",X"70",X"70",X"70",X"70",X"66",
		X"75",X"63",X"1B",X"63",X"1B",X"63",X"23",X"63",X"23",X"63",X"2B",X"63",X"2B",X"63",X"33",X"63",
		X"33",X"63",X"3B",X"63",X"3B",X"63",X"43",X"63",X"43",X"00",X"00",X"72",X"74",X"B6",X"B6",X"B6",
		X"B6",X"B6",X"C7",X"72",X"73",X"74",X"B6",X"B6",X"B6",X"B6",X"C7",X"72",X"73",X"73",X"74",X"B6",
		X"B6",X"B6",X"C7",X"72",X"73",X"73",X"73",X"74",X"B6",X"B6",X"C7",X"72",X"73",X"73",X"73",X"73",
		X"74",X"B6",X"C7",X"72",X"73",X"73",X"73",X"73",X"73",X"74",X"C7",X"BC",X"8B",X"BD",X"8B",X"BE",
		X"8B",X"BF",X"8B",X"AF",X"8A",X"9F",X"89",X"8F",X"88",X"7F",X"87",X"6F",X"86",X"5F",X"85",X"4F",
		X"84",X"3F",X"83",X"2F",X"82",X"1F",X"81",X"0F",X"80",X"0F",X"80",X"6E",X"D8",X"0C",X"FC",X"B8",
		X"92",X"ED",X"49",X"6C",X"48",X"CC",X"63",X"7A",X"ED",X"4C",X"B6",X"B8",X"21",X"26",X"09",X"EC",
		X"49",X"83",X"00",X"01",X"ED",X"49",X"26",X"00",X"10",X"26",X"00",X"8E",X"A6",X"48",X"81",X"06",
		X"25",X"03",X"1A",X"01",X"39",X"31",X"4E",X"CC",X"06",X"02",X"AE",X"22",X"30",X"02",X"AF",X"22",
		X"E7",X"21",X"31",X"24",X"4A",X"26",X"F3",X"CC",X"63",X"B0",X"ED",X"4C",X"6F",X"4B",X"6F",X"49",
		X"6A",X"49",X"2E",X"66",X"86",X"07",X"A7",X"49",X"E6",X"4B",X"CB",X"02",X"E7",X"4B",X"C1",X"10",
		X"22",X"0B",X"8E",X"63",X"49",X"3A",X"EC",X"84",X"FD",X"D0",X"3E",X"20",X"4D",X"CC",X"63",X"D2",
		X"ED",X"4C",X"31",X"4E",X"86",X"06",X"E6",X"21",X"27",X"0C",X"6A",X"21",X"26",X"3C",X"AE",X"22",
		X"30",X"02",X"AF",X"22",X"20",X"34",X"31",X"24",X"4A",X"26",X"EB",X"B6",X"B8",X"29",X"26",X"02",
		X"86",X"0E",X"8B",X"02",X"B7",X"B8",X"29",X"CC",X"63",X"FC",X"ED",X"4C",X"6A",X"49",X"2E",X"1A",
		X"86",X"02",X"A7",X"49",X"E6",X"4B",X"CB",X"FE",X"E7",X"4B",X"2F",X"0B",X"8E",X"63",X"49",X"3A",
		X"EC",X"84",X"FD",X"D0",X"3E",X"20",X"03",X"7E",X"63",X"6E",X"33",X"4E",X"10",X"8E",X"C0",X"51",
		X"CC",X"FF",X"06",X"A7",X"C8",X"14",X"34",X"04",X"8D",X"0C",X"31",X"31",X"33",X"44",X"6A",X"E4",
		X"26",X"F6",X"1C",X"FE",X"35",X"84",X"E6",X"C4",X"5C",X"C1",X"05",X"25",X"01",X"5F",X"E7",X"C4",
		X"AE",X"42",X"AE",X"84",X"58",X"58",X"58",X"3A",X"EC",X"84",X"ED",X"A4",X"EC",X"02",X"ED",X"22",
		X"EC",X"04",X"ED",X"24",X"EC",X"06",X"ED",X"26",X"34",X"20",X"1E",X"20",X"C8",X"F0",X"CB",X"C0",
		X"1E",X"20",X"EC",X"84",X"88",X"80",X"C8",X"80",X"ED",X"A4",X"EC",X"02",X"88",X"80",X"C8",X"80",
		X"ED",X"22",X"EC",X"04",X"88",X"80",X"C8",X"80",X"ED",X"24",X"EC",X"06",X"88",X"80",X"C8",X"80",
		X"ED",X"26",X"35",X"A0",X"CC",X"64",X"8F",X"ED",X"C8",X"5A",X"CC",X"6F",X"C2",X"ED",X"58",X"E6",
		X"5E",X"27",X"55",X"EC",X"5A",X"46",X"56",X"86",X"0A",X"24",X"02",X"8A",X"20",X"97",X"78",X"1F",
		X"98",X"E6",X"5E",X"DD",X"7A",X"AE",X"D8",X"29",X"A3",X"84",X"ED",X"24",X"A3",X"0A",X"ED",X"C8",
		X"52",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"EC",X"08",X"ED",X"44",X"96",X"78",X"A7",
		X"A4",X"31",X"28",X"BD",X"64",X"E9",X"AE",X"C8",X"2B",X"27",X"1A",X"AE",X"84",X"27",X"16",X"DC",
		X"7A",X"A3",X"84",X"ED",X"24",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"96",X"78",X"C6",
		X"88",X"ED",X"A4",X"31",X"28",X"BD",X"65",X"04",X"39",X"A6",X"C8",X"5E",X"2B",X"0A",X"E6",X"C8",
		X"21",X"C5",X"03",X"27",X"03",X"BD",X"65",X"1F",X"AE",X"C8",X"58",X"BC",X"EF",X"D4",X"26",X"03",
		X"7E",X"66",X"0F",X"39",X"A6",X"C8",X"5E",X"2B",X"0A",X"E6",X"C8",X"21",X"C5",X"0C",X"27",X"03",
		X"BD",X"65",X"1F",X"AE",X"C8",X"58",X"BC",X"EF",X"D6",X"26",X"03",X"7E",X"66",X"65",X"39",X"81",
		X"08",X"24",X"39",X"6A",X"C8",X"48",X"2E",X"11",X"86",X"04",X"A7",X"C8",X"48",X"A6",X"C8",X"5E",
		X"8B",X"02",X"A7",X"C8",X"5E",X"81",X"08",X"24",X"20",X"8E",X"66",X"06",X"AB",X"85",X"8E",X"02",
		X"66",X"AE",X"86",X"DC",X"7A",X"A3",X"84",X"ED",X"24",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",
		X"26",X"96",X"78",X"A7",X"A4",X"31",X"28",X"20",X"5B",X"6F",X"C8",X"48",X"6C",X"C8",X"48",X"E6",
		X"C8",X"48",X"C1",X"1E",X"25",X"06",X"86",X"FF",X"A7",X"C8",X"5E",X"39",X"8E",X"02",X"80",X"C4",
		X"06",X"12",X"AE",X"85",X"DC",X"7A",X"A3",X"84",X"ED",X"24",X"EC",X"02",X"ED",X"22",X"EC",X"06",
		X"ED",X"26",X"96",X"78",X"A7",X"A4",X"E6",X"C8",X"48",X"54",X"E1",X"27",X"24",X"13",X"A6",X"27",
		X"E7",X"27",X"A0",X"27",X"1F",X"89",X"AB",X"25",X"A7",X"25",X"A6",X"26",X"3D",X"E3",X"22",X"ED",
		X"22",X"8E",X"65",X"F3",X"A6",X"C8",X"21",X"E6",X"86",X"8E",X"65",X"FC",X"EC",X"85",X"E3",X"24",
		X"ED",X"24",X"31",X"28",X"A6",X"C8",X"52",X"A0",X"3C",X"23",X"09",X"AB",X"44",X"A7",X"44",X"A6",
		X"3C",X"A7",X"C8",X"52",X"A6",X"3C",X"AB",X"3E",X"A0",X"C8",X"52",X"A0",X"44",X"2F",X"04",X"AB",
		X"44",X"A7",X"44",X"E6",X"C8",X"53",X"E0",X"3D",X"23",X"09",X"EB",X"45",X"E7",X"45",X"E6",X"3D",
		X"E7",X"C8",X"53",X"E6",X"3D",X"EB",X"3F",X"E0",X"C8",X"53",X"E0",X"45",X"2F",X"04",X"EB",X"45",
		X"E7",X"45",X"39",X"00",X"02",X"04",X"00",X"06",X"00",X"00",X"00",X"08",X"00",X"00",X"03",X"FA",
		X"FB",X"FA",X"04",X"06",X"FC",X"06",X"00",X"00",X"06",X"00",X"0C",X"00",X"00",X"00",X"12",X"6A",
		X"C8",X"18",X"2E",X"24",X"86",X"04",X"A7",X"C8",X"18",X"6C",X"C8",X"19",X"A6",X"C8",X"19",X"81",
		X"05",X"22",X"5B",X"81",X"03",X"26",X"11",X"5F",X"A6",X"C8",X"20",X"85",X"09",X"26",X"02",X"CB",
		X"0A",X"8E",X"02",X"46",X"3A",X"AF",X"C8",X"29",X"8E",X"02",X"98",X"A6",X"C8",X"20",X"85",X"0A",
		X"27",X"02",X"30",X"08",X"E6",X"C8",X"19",X"58",X"3A",X"AE",X"84",X"DC",X"7A",X"A3",X"84",X"ED",
		X"24",X"ED",X"C8",X"5C",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"ED",X"46",X"96",X"78",
		X"A7",X"A4",X"31",X"28",X"39",X"6A",X"C8",X"18",X"2E",X"1E",X"5F",X"4F",X"ED",X"C8",X"2B",X"86",
		X"04",X"A7",X"C8",X"18",X"6C",X"C8",X"19",X"A6",X"C8",X"19",X"81",X"05",X"23",X"0A",X"CC",X"6F",
		X"EA",X"ED",X"C8",X"58",X"6F",X"C8",X"18",X"39",X"8E",X"02",X"88",X"A6",X"C8",X"21",X"20",X"AE",
		X"3F",X"39",X"CC",X"66",X"A0",X"ED",X"C8",X"5A",X"CC",X"6F",X"C2",X"ED",X"58",X"6F",X"C8",X"33",
		X"E6",X"5E",X"26",X"01",X"39",X"EC",X"5A",X"46",X"56",X"86",X"0A",X"24",X"02",X"8A",X"20",X"97",
		X"78",X"1F",X"98",X"E6",X"5E",X"DD",X"7A",X"A6",X"C8",X"39",X"81",X"10",X"24",X"6E",X"1F",X"89",
		X"34",X"06",X"8E",X"02",X"F6",X"6C",X"C8",X"33",X"E6",X"C8",X"33",X"C4",X"03",X"58",X"AE",X"85",
		X"DC",X"7A",X"A3",X"84",X"ED",X"24",X"A3",X"0A",X"ED",X"C8",X"52",X"EC",X"02",X"ED",X"22",X"A6",
		X"06",X"E6",X"61",X"CB",X"04",X"E1",X"07",X"25",X"02",X"E6",X"07",X"ED",X"26",X"EC",X"08",X"ED",
		X"44",X"E6",X"07",X"E0",X"27",X"1F",X"98",X"E7",X"E4",X"EB",X"25",X"E7",X"25",X"E6",X"26",X"3D",
		X"E3",X"22",X"ED",X"22",X"96",X"78",X"A7",X"A4",X"31",X"28",X"BE",X"02",X"FE",X"DC",X"7A",X"A3",
		X"84",X"60",X"61",X"EB",X"61",X"ED",X"24",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"96",
		X"78",X"8A",X"10",X"E6",X"C8",X"37",X"ED",X"A4",X"31",X"28",X"35",X"86",X"1F",X"89",X"C1",X"1C",
		X"22",X"0A",X"50",X"CB",X"1F",X"C1",X"08",X"2D",X"03",X"7E",X"66",X"C0",X"A6",X"C8",X"35",X"26",
		X"03",X"6C",X"C8",X"35",X"AE",X"D8",X"29",X"DC",X"7A",X"A3",X"84",X"A3",X"0A",X"ED",X"C8",X"52",
		X"EC",X"08",X"ED",X"44",X"AE",X"D8",X"29",X"DC",X"7A",X"A3",X"84",X"ED",X"24",X"A3",X"0A",X"34",
		X"06",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"96",X"78",X"A7",X"A4",X"31",X"28",X"C6",
		X"0B",X"A6",X"C8",X"39",X"3D",X"40",X"8B",X"08",X"2A",X"01",X"4F",X"1F",X"89",X"BD",X"66",X"C0",
		X"35",X"06",X"ED",X"C8",X"52",X"AE",X"D8",X"29",X"EC",X"08",X"ED",X"44",X"AE",X"D8",X"2B",X"DC",
		X"7A",X"A3",X"84",X"ED",X"24",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"96",X"78",X"A7",
		X"A4",X"31",X"28",X"39",X"CC",X"67",X"AF",X"ED",X"C8",X"5A",X"CC",X"6F",X"C2",X"ED",X"58",X"E6",
		X"5E",X"26",X"01",X"39",X"EC",X"5A",X"46",X"56",X"86",X"0A",X"24",X"02",X"8A",X"20",X"97",X"78",
		X"1F",X"98",X"E6",X"5E",X"DD",X"7A",X"0F",X"79",X"A6",X"C8",X"21",X"26",X"0A",X"A6",X"C8",X"10",
		X"E6",X"C8",X"3B",X"10",X"27",X"00",X"9E",X"85",X"0C",X"27",X"04",X"C6",X"07",X"D7",X"79",X"EC",
		X"C8",X"18",X"E3",X"C8",X"14",X"1F",X"01",X"A6",X"89",X"91",X"02",X"2B",X"0F",X"85",X"0F",X"27",
		X"0B",X"E6",X"C8",X"48",X"C4",X"06",X"26",X"0E",X"85",X"10",X"26",X"0A",X"E6",X"C8",X"10",X"8E",
		X"68",X"B2",X"E6",X"85",X"20",X"23",X"CB",X"FE",X"2A",X"02",X"CB",X"06",X"A6",X"C8",X"10",X"85",
		X"03",X"27",X"08",X"CB",X"04",X"C1",X"06",X"2D",X"02",X"C0",X"06",X"58",X"58",X"58",X"EB",X"C8",
		X"48",X"CA",X"08",X"85",X"09",X"27",X"02",X"C4",X"F7",X"D7",X"7F",X"8E",X"01",X"CC",X"3A",X"3A",
		X"EC",X"02",X"D3",X"7A",X"AE",X"84",X"A3",X"84",X"DD",X"7D",X"EB",X"0C",X"ED",X"24",X"EC",X"02",
		X"ED",X"22",X"EC",X"06",X"ED",X"26",X"96",X"78",X"ED",X"A4",X"31",X"28",X"D6",X"7F",X"CA",X"08",
		X"C1",X"2A",X"26",X"21",X"D6",X"7F",X"C4",X"08",X"CB",X"26",X"8E",X"01",X"CC",X"3A",X"3A",X"EC",
		X"02",X"D3",X"7D",X"AE",X"84",X"ED",X"24",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"96",
		X"78",X"ED",X"A4",X"31",X"28",X"AE",X"D8",X"29",X"DC",X"7A",X"A3",X"84",X"ED",X"24",X"A3",X"0A",
		X"ED",X"C8",X"52",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"EC",X"08",X"DB",X"79",X"ED",
		X"44",X"96",X"78",X"A7",X"A4",X"31",X"28",X"AE",X"D8",X"2B",X"DC",X"7A",X"A3",X"84",X"ED",X"24",
		X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"96",X"78",X"A7",X"A4",X"31",X"28",X"AD",X"D8",
		X"58",X"39",X"00",X"06",X"0E",X"00",X"16",X"00",X"00",X"00",X"1E",X"CC",X"68",X"D1",X"ED",X"C8",
		X"5A",X"CC",X"F8",X"00",X"ED",X"C8",X"35",X"4F",X"5F",X"ED",X"C8",X"33",X"CC",X"6A",X"53",X"ED",
		X"58",X"EC",X"5D",X"26",X"01",X"39",X"EC",X"5A",X"46",X"56",X"86",X"0A",X"24",X"02",X"8A",X"20",
		X"97",X"78",X"1F",X"98",X"E6",X"5E",X"DD",X"7A",X"AE",X"D8",X"29",X"27",X"2A",X"A6",X"C8",X"18",
		X"81",X"04",X"22",X"23",X"34",X"01",X"DC",X"7A",X"A3",X"84",X"ED",X"24",X"EC",X"06",X"ED",X"26",
		X"EC",X"02",X"ED",X"22",X"96",X"78",X"5F",X"35",X"01",X"26",X"08",X"E7",X"C8",X"29",X"E7",X"C8",
		X"2A",X"8A",X"10",X"ED",X"A4",X"31",X"28",X"6A",X"C8",X"19",X"2E",X"0D",X"86",X"04",X"A7",X"C8",
		X"19",X"6C",X"C8",X"18",X"2E",X"03",X"6A",X"C8",X"18",X"8E",X"02",X"C2",X"A6",X"C8",X"18",X"81",
		X"05",X"22",X"1C",X"48",X"AE",X"86",X"DC",X"7A",X"A3",X"84",X"ED",X"24",X"ED",X"C8",X"52",X"EC",
		X"06",X"ED",X"26",X"ED",X"44",X"EC",X"02",X"ED",X"22",X"96",X"78",X"A7",X"A4",X"31",X"28",X"CC",
		X"00",X"40",X"E3",X"C8",X"35",X"10",X"83",X"08",X"00",X"2E",X"03",X"ED",X"C8",X"35",X"A6",X"C8",
		X"10",X"48",X"8E",X"69",X"AA",X"EC",X"86",X"E3",X"C8",X"33",X"EB",X"C8",X"35",X"ED",X"C8",X"33",
		X"AE",X"D8",X"2B",X"DC",X"7A",X"A3",X"84",X"AB",X"C8",X"33",X"81",X"90",X"22",X"1D",X"EB",X"C8",
		X"34",X"C1",X"F0",X"22",X"16",X"ED",X"24",X"ED",X"C8",X"5C",X"EC",X"06",X"ED",X"26",X"ED",X"46",
		X"EC",X"02",X"ED",X"22",X"96",X"78",X"A7",X"A4",X"31",X"28",X"39",X"A6",X"C8",X"18",X"81",X"05",
		X"25",X"09",X"6F",X"C8",X"18",X"CC",X"6F",X"EA",X"ED",X"C8",X"5A",X"39",X"01",X"03",X"FF",X"03",
		X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",X"CC",X"69",X"C7",X"ED",
		X"C8",X"5A",X"CC",X"6A",X"53",X"ED",X"58",X"EC",X"5D",X"26",X"01",X"39",X"EC",X"5A",X"46",X"56",
		X"86",X"0A",X"24",X"02",X"8A",X"20",X"97",X"78",X"1F",X"98",X"E6",X"5E",X"DD",X"7A",X"C6",X"FF",
		X"E7",X"C8",X"43",X"AE",X"C8",X"14",X"8C",X"09",X"40",X"24",X"30",X"E6",X"89",X"91",X"02",X"2B",
		X"2A",X"C5",X"0F",X"27",X"26",X"54",X"54",X"C4",X"3C",X"50",X"EB",X"42",X"DB",X"7B",X"AE",X"D8",
		X"29",X"AE",X"04",X"A3",X"84",X"ED",X"24",X"ED",X"C8",X"41",X"EC",X"02",X"ED",X"22",X"EC",X"06",
		X"ED",X"26",X"ED",X"C8",X"43",X"96",X"78",X"A7",X"A4",X"31",X"28",X"AE",X"D8",X"29",X"DC",X"7A",
		X"A3",X"84",X"ED",X"24",X"A3",X"0A",X"ED",X"C8",X"52",X"EC",X"06",X"ED",X"26",X"EC",X"02",X"ED",
		X"22",X"EC",X"08",X"ED",X"44",X"96",X"78",X"A7",X"A4",X"31",X"28",X"AE",X"D8",X"2B",X"DC",X"7A",
		X"A3",X"84",X"ED",X"24",X"EC",X"06",X"ED",X"26",X"EC",X"02",X"ED",X"22",X"96",X"78",X"A7",X"A4",
		X"31",X"28",X"39",X"EC",X"44",X"2F",X"23",X"60",X"44",X"ED",X"26",X"EC",X"C8",X"52",X"ED",X"24",
		X"CC",X"12",X"00",X"ED",X"A4",X"31",X"28",X"ED",X"A4",X"EC",X"C8",X"43",X"2F",X"0C",X"60",X"C8",
		X"43",X"ED",X"26",X"EC",X"C8",X"41",X"ED",X"24",X"31",X"28",X"EC",X"46",X"2F",X"10",X"60",X"46",
		X"ED",X"26",X"EC",X"C8",X"5C",X"ED",X"24",X"CC",X"12",X"00",X"ED",X"A4",X"31",X"28",X"39",X"CC",
		X"6A",X"9A",X"ED",X"C8",X"5A",X"CC",X"6B",X"09",X"ED",X"58",X"E6",X"5E",X"27",X"6A",X"CC",X"00",
		X"00",X"ED",X"C8",X"52",X"EC",X"5A",X"46",X"56",X"86",X"0A",X"24",X"02",X"8A",X"20",X"97",X"78",
		X"1F",X"98",X"E6",X"5E",X"DD",X"7A",X"AE",X"C8",X"14",X"E6",X"89",X"91",X"02",X"2B",X"2D",X"C5",
		X"0F",X"27",X"29",X"54",X"54",X"C4",X"3C",X"50",X"EB",X"42",X"EB",X"5E",X"CB",X"00",X"AE",X"D8",
		X"2D",X"A3",X"84",X"ED",X"24",X"ED",X"C8",X"5C",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",
		X"ED",X"46",X"96",X"78",X"8A",X"10",X"C6",X"88",X"ED",X"A4",X"31",X"28",X"AE",X"D8",X"29",X"DC",
		X"7A",X"A3",X"84",X"ED",X"24",X"ED",X"C8",X"52",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",
		X"ED",X"44",X"96",X"78",X"A7",X"A4",X"31",X"28",X"39",X"EC",X"44",X"2F",X"10",X"60",X"44",X"ED",
		X"26",X"EC",X"C8",X"52",X"ED",X"24",X"CC",X"12",X"00",X"ED",X"A4",X"31",X"28",X"EC",X"46",X"2F",
		X"10",X"60",X"46",X"ED",X"26",X"EC",X"C8",X"5C",X"ED",X"24",X"CC",X"12",X"00",X"ED",X"A4",X"31",
		X"28",X"39",X"CC",X"6B",X"3D",X"ED",X"C8",X"5A",X"CC",X"6B",X"B0",X"ED",X"58",X"E6",X"5E",X"27",
		X"6E",X"CC",X"00",X"00",X"ED",X"C8",X"52",X"EC",X"5A",X"46",X"56",X"86",X"0A",X"24",X"02",X"8A",
		X"20",X"97",X"78",X"1F",X"98",X"E6",X"5E",X"DD",X"7A",X"AE",X"C8",X"14",X"8C",X"09",X"40",X"24",
		X"32",X"E6",X"89",X"91",X"02",X"2B",X"2C",X"C5",X"0F",X"27",X"28",X"54",X"54",X"C4",X"3C",X"50",
		X"EB",X"C8",X"5E",X"2F",X"1E",X"EB",X"5E",X"AE",X"D8",X"29",X"A3",X"84",X"ED",X"24",X"ED",X"C8",
		X"52",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"96",X"78",X"8A",X"10",X"C6",X"88",X"ED",
		X"A4",X"31",X"28",X"AE",X"D8",X"29",X"DC",X"7A",X"A3",X"84",X"ED",X"24",X"ED",X"C8",X"4B",X"EC",
		X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"ED",X"44",X"96",X"78",X"A7",X"A4",X"31",X"28",X"39",
		X"EC",X"44",X"2F",X"1A",X"60",X"44",X"ED",X"26",X"ED",X"2E",X"EC",X"C8",X"4B",X"ED",X"24",X"EC",
		X"C8",X"52",X"ED",X"2C",X"CC",X"12",X"00",X"ED",X"A4",X"ED",X"28",X"31",X"A8",X"10",X"EC",X"46",
		X"2F",X"10",X"60",X"46",X"ED",X"26",X"EC",X"C8",X"5C",X"ED",X"24",X"CC",X"12",X"00",X"ED",X"A4",
		X"31",X"28",X"39",X"CC",X"6B",X"EE",X"ED",X"C8",X"5A",X"CC",X"6F",X"C2",X"ED",X"58",X"E6",X"5E",
		X"27",X"2E",X"EC",X"5A",X"46",X"56",X"86",X"0A",X"24",X"02",X"8A",X"20",X"97",X"78",X"1F",X"98",
		X"E6",X"5E",X"DD",X"7A",X"AE",X"D8",X"29",X"DC",X"7A",X"A3",X"84",X"ED",X"24",X"ED",X"C8",X"52",
		X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"ED",X"44",X"96",X"78",X"A7",X"A4",X"31",X"28",
		X"39",X"CC",X"6C",X"2C",X"ED",X"C8",X"58",X"86",X"0C",X"A7",X"C8",X"5C",X"6A",X"C8",X"5C",X"2F",
		X"2A",X"8E",X"6C",X"4B",X"E6",X"C8",X"5C",X"3A",X"EC",X"30",X"E6",X"84",X"27",X"0C",X"8A",X"10",
		X"ED",X"30",X"EC",X"38",X"E6",X"84",X"8A",X"10",X"ED",X"38",X"39",X"EE",X"00",X"EE",X"00",X"11",
		X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"6F",X"C8",X"5C",X"CC",X"6C",
		X"64",X"ED",X"C8",X"58",X"39",X"CC",X"6C",X"70",X"ED",X"C8",X"58",X"86",X"10",X"A7",X"C8",X"5C",
		X"6A",X"C8",X"5C",X"2B",X"2F",X"8E",X"6C",X"94",X"E6",X"C8",X"5C",X"3A",X"E6",X"84",X"27",X"13",
		X"C1",X"01",X"26",X"03",X"E6",X"C8",X"5D",X"A6",X"30",X"8A",X"10",X"ED",X"30",X"A6",X"38",X"8A",
		X"10",X"ED",X"38",X"39",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"01",X"00",X"01",
		X"01",X"00",X"01",X"01",X"CC",X"6C",X"AA",X"ED",X"C8",X"58",X"39",X"CC",X"6F",X"C2",X"ED",X"58",
		X"EC",X"5A",X"46",X"56",X"86",X"0A",X"24",X"02",X"8A",X"20",X"97",X"78",X"1F",X"98",X"E6",X"5E",
		X"DD",X"7A",X"8E",X"B2",X"EE",X"A6",X"51",X"81",X"01",X"27",X"03",X"8E",X"B5",X"02",X"AF",X"C8",
		X"42",X"34",X"01",X"1A",X"F0",X"BD",X"6E",X"4F",X"AE",X"D8",X"29",X"CC",X"07",X"FF",X"A3",X"84",
		X"FD",X"C8",X"84",X"A3",X"0A",X"ED",X"C8",X"52",X"EC",X"02",X"FD",X"C8",X"82",X"EC",X"06",X"FD",
		X"C8",X"86",X"EC",X"08",X"ED",X"44",X"ED",X"C8",X"40",X"96",X"78",X"BD",X"E0",X"96",X"AE",X"D8",
		X"2B",X"CC",X"07",X"FF",X"A3",X"84",X"FD",X"C8",X"84",X"EC",X"02",X"FD",X"C8",X"82",X"EC",X"06",
		X"FD",X"C8",X"86",X"96",X"78",X"BD",X"E0",X"96",X"AE",X"C8",X"42",X"BF",X"C8",X"84",X"EC",X"C8",
		X"52",X"FD",X"C8",X"82",X"EC",X"44",X"FD",X"C8",X"86",X"86",X"05",X"BD",X"E0",X"90",X"BD",X"6E",
		X"4F",X"35",X"01",X"AE",X"D8",X"29",X"DC",X"7A",X"A3",X"84",X"A3",X"0A",X"ED",X"C8",X"52",X"ED",
		X"C8",X"46",X"86",X"20",X"A7",X"C8",X"3E",X"39",X"CC",X"6D",X"5A",X"ED",X"C8",X"5A",X"BD",X"6C",
		X"AB",X"A6",X"C8",X"40",X"4C",X"48",X"48",X"A7",X"C8",X"3E",X"E6",X"5E",X"26",X"01",X"39",X"AE",
		X"C8",X"42",X"AF",X"22",X"EC",X"C8",X"40",X"ED",X"44",X"ED",X"26",X"EC",X"C8",X"46",X"ED",X"C8",
		X"52",X"ED",X"24",X"86",X"0E",X"A7",X"A4",X"31",X"28",X"A6",X"C8",X"3E",X"84",X"03",X"26",X"36",
		X"EC",X"3E",X"4C",X"44",X"34",X"16",X"86",X"04",X"1C",X"FE",X"AE",X"62",X"E6",X"E4",X"66",X"80",
		X"5A",X"26",X"FB",X"4A",X"26",X"F2",X"86",X"04",X"1C",X"FE",X"AE",X"62",X"E6",X"3E",X"3A",X"E6",
		X"E4",X"69",X"82",X"5A",X"26",X"FB",X"4A",X"26",X"EF",X"AE",X"62",X"E6",X"3E",X"3A",X"AF",X"62",
		X"6A",X"61",X"26",X"D2",X"35",X"16",X"39",X"CC",X"6D",X"C0",X"ED",X"C8",X"5A",X"BD",X"6C",X"AB",
		X"E6",X"5E",X"26",X"01",X"39",X"AE",X"C8",X"42",X"AF",X"22",X"EC",X"C8",X"40",X"ED",X"44",X"ED",
		X"26",X"EC",X"C8",X"46",X"ED",X"C8",X"52",X"ED",X"24",X"86",X"0E",X"A7",X"A4",X"31",X"28",X"A6",
		X"C8",X"3E",X"44",X"25",X"04",X"85",X"01",X"26",X"08",X"A6",X"38",X"C6",X"99",X"8A",X"10",X"ED",
		X"38",X"A6",X"C8",X"3E",X"44",X"24",X"17",X"E6",X"C8",X"3E",X"C4",X"06",X"8E",X"6E",X"47",X"3A",
		X"EC",X"84",X"E3",X"3C",X"ED",X"3C",X"EC",X"84",X"E3",X"C8",X"52",X"ED",X"C8",X"52",X"E6",X"C8",
		X"40",X"86",X"20",X"A0",X"C8",X"3E",X"3D",X"E3",X"C8",X"42",X"1F",X"01",X"E6",X"C8",X"40",X"5A",
		X"54",X"D7",X"7A",X"E6",X"C8",X"40",X"50",X"1D",X"DD",X"78",X"4F",X"E6",X"C8",X"40",X"5A",X"6F",
		X"86",X"6F",X"85",X"4C",X"5A",X"91",X"7A",X"22",X"0D",X"1E",X"10",X"D3",X"78",X"D3",X"78",X"1E",
		X"01",X"AC",X"C8",X"42",X"24",X"E9",X"39",X"FF",X"FE",X"01",X"00",X"00",X"02",X"FF",X"00",X"CC",
		X"0E",X"2A",X"FD",X"C8",X"86",X"CC",X"00",X"D5",X"FD",X"C8",X"84",X"CC",X"12",X"00",X"F7",X"C8",
		X"81",X"B7",X"C8",X"80",X"39",X"CC",X"6E",X"70",X"ED",X"C8",X"5A",X"CC",X"6F",X"C2",X"ED",X"58",
		X"E6",X"5E",X"27",X"66",X"AE",X"D8",X"29",X"EC",X"5A",X"46",X"56",X"86",X"0A",X"24",X"02",X"8A",
		X"20",X"7D",X"B7",X"48",X"26",X"05",X"6D",X"C8",X"51",X"2A",X"02",X"8A",X"10",X"97",X"78",X"1F",
		X"98",X"E6",X"5E",X"DD",X"7A",X"EB",X"C8",X"5E",X"A3",X"84",X"ED",X"24",X"E0",X"0B",X"A0",X"0A",
		X"ED",X"C8",X"52",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"EC",X"08",X"ED",X"44",X"96",
		X"78",X"C6",X"88",X"ED",X"A4",X"31",X"28",X"A6",X"C8",X"5E",X"81",X"F4",X"2F",X"1C",X"AE",X"D8",
		X"2B",X"DC",X"7A",X"A3",X"84",X"ED",X"24",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"96",
		X"78",X"C6",X"88",X"ED",X"A4",X"31",X"28",X"AD",X"D8",X"58",X"39",X"CC",X"6E",X"E6",X"ED",X"C8",
		X"5A",X"CC",X"6F",X"C2",X"ED",X"58",X"B6",X"B8",X"31",X"27",X"62",X"E6",X"5E",X"27",X"5D",X"AE",
		X"D8",X"29",X"EC",X"5A",X"46",X"56",X"86",X"0A",X"24",X"02",X"8A",X"20",X"97",X"78",X"1F",X"98",
		X"E6",X"5E",X"DD",X"7A",X"A3",X"84",X"ED",X"24",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",
		X"96",X"78",X"A7",X"A4",X"31",X"28",X"AE",X"D8",X"2B",X"DC",X"7A",X"A3",X"84",X"ED",X"24",X"EC",
		X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"96",X"78",X"A7",X"A4",X"31",X"28",X"BE",X"03",X"24",
		X"DC",X"7A",X"A3",X"84",X"ED",X"24",X"ED",X"C8",X"52",X"CC",X"BE",X"1F",X"ED",X"22",X"EC",X"06",
		X"ED",X"26",X"ED",X"44",X"96",X"78",X"8A",X"04",X"A7",X"A4",X"31",X"28",X"39",X"CC",X"6F",X"58",
		X"ED",X"C8",X"5A",X"CC",X"6F",X"C2",X"ED",X"58",X"E6",X"5E",X"27",X"65",X"AE",X"D8",X"29",X"EC",
		X"5A",X"46",X"56",X"86",X"0A",X"24",X"02",X"8A",X"20",X"7D",X"B7",X"48",X"26",X"05",X"6D",X"C8",
		X"51",X"2A",X"02",X"8A",X"10",X"97",X"78",X"1F",X"98",X"E6",X"5E",X"DD",X"7A",X"A3",X"84",X"ED",
		X"24",X"A3",X"0A",X"ED",X"C8",X"52",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"EC",X"08",
		X"ED",X"44",X"96",X"78",X"C6",X"88",X"ED",X"A4",X"31",X"28",X"AE",X"C8",X"2B",X"96",X"78",X"C6",
		X"88",X"7D",X"B7",X"48",X"27",X"04",X"30",X"08",X"84",X"EF",X"ED",X"A4",X"AE",X"84",X"DC",X"7A",
		X"A3",X"84",X"ED",X"24",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"31",X"28",X"AD",X"D8",
		X"58",X"39",X"EC",X"44",X"2F",X"10",X"60",X"44",X"ED",X"26",X"EC",X"C8",X"52",X"ED",X"24",X"CC",
		X"12",X"00",X"ED",X"A4",X"31",X"28",X"EC",X"46",X"2F",X"10",X"60",X"46",X"ED",X"26",X"EC",X"C8",
		X"5C",X"ED",X"24",X"CC",X"12",X"00",X"ED",X"A4",X"31",X"28",X"39",X"3F",X"39",X"20",X"49",X"4E",
		X"46",X"45",X"52",X"4E",X"4F",X"20",X"2D",X"20",X"28",X"43",X"29",X"31",X"39",X"38",X"34",X"20",
		X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",
		X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
