library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity inferno_graph2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of inferno_graph2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"02",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"00",X"11",X"11",X"00",X"02",X"11",X"12",X"00",X"11",X"11",X"37",X"00",X"11",X"11",X"09",
		X"00",X"11",X"11",X"00",X"02",X"11",X"12",X"00",X"11",X"11",X"39",X"00",X"11",X"11",X"09",X"00",
		X"11",X"11",X"08",X"00",X"11",X"12",X"00",X"00",X"11",X"37",X"00",X"00",X"11",X"09",X"00",X"00",
		X"11",X"09",X"00",X"00",X"12",X"08",X"00",X"00",X"39",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"37",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"00",X"00",X"72",X"12",X"00",X"00",X"07",X"37",X"00",X"00",X"09",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"00",X"00",X"00",X"12",X"00",X"00",X"02",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",
		X"11",X"30",X"00",X"11",X"11",X"12",X"02",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"92",X"11",X"11",X"12",X"97",X"11",X"11",X"37",X"80",X"11",X"11",X"09",
		X"00",X"11",X"11",X"00",X"02",X"11",X"12",X"00",X"11",X"11",X"37",X"00",X"11",X"11",X"09",X"00",
		X"11",X"11",X"09",X"00",X"11",X"12",X"08",X"00",X"11",X"39",X"00",X"00",X"11",X"09",X"00",X"00",
		X"11",X"38",X"00",X"00",X"11",X"12",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",
		X"11",X"11",X"30",X"00",X"72",X"11",X"12",X"00",X"07",X"11",X"11",X"00",X"09",X"11",X"11",X"00",
		X"00",X"11",X"11",X"30",X"02",X"11",X"11",X"12",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"12",X"72",X"11",X"11",X"39",X"07",X"11",X"11",X"09",X"09",X"11",
		X"11",X"08",X"00",X"11",X"12",X"00",X"00",X"72",X"37",X"00",X"00",X"07",X"09",X"00",X"00",X"09",
		X"09",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"00",X"02",X"11",X"12",X"00",X"11",X"11",X"39",X"00",X"11",X"11",X"09",X"00",
		X"11",X"11",X"08",X"00",X"11",X"12",X"00",X"02",X"11",X"37",X"00",X"11",X"11",X"09",X"00",X"11",
		X"11",X"09",X"00",X"11",X"12",X"08",X"02",X"11",X"39",X"00",X"11",X"11",X"09",X"00",X"11",X"11",
		X"08",X"00",X"11",X"11",X"00",X"02",X"11",X"12",X"00",X"11",X"11",X"37",X"00",X"11",X"11",X"09",
		X"00",X"11",X"11",X"30",X"00",X"72",X"11",X"12",X"00",X"07",X"11",X"11",X"00",X"09",X"11",X"11",
		X"30",X"00",X"11",X"11",X"12",X"00",X"72",X"11",X"11",X"00",X"07",X"11",X"11",X"00",X"09",X"11",
		X"11",X"30",X"00",X"11",X"11",X"12",X"02",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"72",X"11",X"11",X"12",X"07",X"11",X"11",X"37",X"09",X"11",X"11",X"09",
		X"00",X"11",X"11",X"30",X"02",X"11",X"11",X"12",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"12",X"72",X"11",X"11",X"37",X"07",X"11",X"11",X"09",X"09",X"11",
		X"11",X"30",X"00",X"11",X"11",X"12",X"00",X"72",X"11",X"11",X"00",X"07",X"11",X"11",X"00",X"09",
		X"11",X"11",X"30",X"00",X"72",X"11",X"12",X"00",X"07",X"11",X"11",X"00",X"09",X"11",X"11",X"00",
		X"00",X"11",X"11",X"30",X"02",X"11",X"11",X"12",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"12",X"72",X"11",X"11",X"37",X"07",X"11",X"11",X"00",X"09",X"11",
		X"11",X"30",X"00",X"11",X"11",X"12",X"02",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"72",X"11",X"11",X"12",X"07",X"11",X"11",X"39",X"09",X"11",X"11",X"09",
		X"00",X"11",X"11",X"00",X"00",X"72",X"12",X"00",X"00",X"07",X"37",X"00",X"00",X"09",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"08",X"02",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"02",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"00",X"11",X"11",X"00",X"02",X"11",X"12",X"00",X"11",X"11",X"37",X"00",X"11",X"11",X"09",
		X"00",X"11",X"11",X"00",X"00",X"21",X"11",X"20",X"00",X"93",X"11",X"11",X"00",X"90",X"11",X"11",
		X"00",X"80",X"11",X"11",X"00",X"00",X"21",X"11",X"00",X"00",X"73",X"11",X"00",X"00",X"90",X"11",
		X"00",X"00",X"90",X"11",X"00",X"00",X"80",X"21",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"90",
		X"00",X"00",X"30",X"80",X"00",X"02",X"12",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",
		X"00",X"11",X"11",X"00",X"00",X"72",X"12",X"00",X"00",X"07",X"37",X"00",X"00",X"09",X"09",X"00",
		X"00",X"00",X"09",X"03",X"00",X"00",X"08",X"21",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"73",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"00",X"00",X"72",X"12",X"00",X"00",X"07",X"37",X"00",X"00",X"09",X"09",X"00",
		X"30",X"00",X"09",X"00",X"12",X"00",X"08",X"02",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",
		X"11",X"30",X"00",X"11",X"11",X"12",X"02",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"92",X"11",X"11",X"12",X"97",X"11",X"11",X"37",X"80",X"11",X"11",X"09",
		X"00",X"11",X"11",X"00",X"00",X"21",X"11",X"20",X"00",X"73",X"11",X"11",X"00",X"90",X"11",X"11",
		X"30",X"90",X"11",X"11",X"12",X"80",X"21",X"11",X"11",X"00",X"93",X"11",X"11",X"00",X"90",X"11",
		X"11",X"00",X"83",X"11",X"12",X"00",X"21",X"11",X"37",X"00",X"11",X"11",X"09",X"00",X"11",X"11",
		X"09",X"03",X"11",X"11",X"08",X"21",X"11",X"27",X"00",X"11",X"11",X"70",X"00",X"11",X"11",X"90",
		X"00",X"11",X"11",X"30",X"02",X"11",X"11",X"12",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"12",X"72",X"11",X"11",X"39",X"07",X"11",X"11",X"09",X"09",X"11",
		X"11",X"08",X"00",X"11",X"12",X"00",X"00",X"72",X"37",X"00",X"00",X"07",X"09",X"00",X"00",X"09",
		X"09",X"00",X"30",X"00",X"08",X"02",X"12",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",
		X"44",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"67",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"08",X"00",X"00",X"02",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"02",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"00",X"11",X"11",X"00",X"02",X"11",X"12",X"00",X"11",X"11",X"37",X"00",X"11",X"11",X"09",
		X"00",X"11",X"11",X"00",X"00",X"21",X"11",X"20",X"00",X"93",X"11",X"11",X"00",X"90",X"11",X"11",
		X"00",X"80",X"11",X"11",X"00",X"00",X"21",X"11",X"00",X"00",X"73",X"11",X"00",X"00",X"90",X"11",
		X"00",X"00",X"90",X"11",X"00",X"00",X"80",X"21",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"80",X"50",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"67",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"03",X"08",X"00",X"00",X"21",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"73",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"67",X"00",X"00",X"00",X"77",X"12",X"00",X"00",
		X"77",X"37",X"00",X"00",X"72",X"77",X"00",X"02",X"11",X"77",X"00",X"11",X"12",X"72",X"00",X"11",
		X"97",X"11",X"00",X"11",X"07",X"12",X"02",X"11",X"07",X"37",X"11",X"11",X"02",X"77",X"11",X"11",
		X"07",X"77",X"11",X"11",X"09",X"72",X"11",X"12",X"09",X"11",X"11",X"37",X"08",X"11",X"11",X"00",
		X"00",X"11",X"11",X"00",X"02",X"11",X"12",X"00",X"11",X"11",X"37",X"00",X"11",X"11",X"77",X"45",
		X"11",X"11",X"77",X"67",X"11",X"12",X"75",X"77",X"11",X"37",X"44",X"77",X"11",X"09",X"45",X"75",
		X"11",X"09",X"97",X"44",X"12",X"08",X"07",X"45",X"39",X"00",X"07",X"67",X"09",X"00",X"05",X"77",
		X"08",X"00",X"07",X"77",X"00",X"00",X"09",X"75",X"00",X"00",X"09",X"44",X"00",X"00",X"08",X"44",
		X"44",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"67",X"00",X"00",X"00",X"77",X"12",X"00",X"00",
		X"77",X"37",X"00",X"00",X"72",X"77",X"00",X"00",X"11",X"77",X"00",X"00",X"12",X"72",X"00",X"00",
		X"97",X"11",X"00",X"00",X"07",X"12",X"00",X"00",X"07",X"37",X"00",X"00",X"02",X"77",X"00",X"00",
		X"07",X"77",X"30",X"00",X"09",X"72",X"12",X"00",X"09",X"11",X"11",X"00",X"08",X"11",X"11",X"00",
		X"00",X"11",X"11",X"00",X"00",X"72",X"12",X"00",X"00",X"07",X"37",X"00",X"00",X"09",X"77",X"45",
		X"00",X"00",X"77",X"67",X"00",X"00",X"75",X"77",X"00",X"00",X"44",X"77",X"00",X"00",X"45",X"75",
		X"00",X"00",X"97",X"44",X"00",X"00",X"07",X"45",X"00",X"00",X"07",X"67",X"00",X"00",X"05",X"77",
		X"00",X"00",X"07",X"77",X"00",X"00",X"09",X"75",X"00",X"00",X"09",X"44",X"00",X"00",X"08",X"44",
		X"00",X"0E",X"2B",X"00",X"C4",X"EB",X"B2",X"00",X"44",X"BC",X"0B",X"B0",X"44",X"C1",X"90",X"2B",
		X"04",X"A1",X"11",X"22",X"DB",X"AA",X"10",X"23",X"0B",X"AA",X"2C",X"33",X"DD",X"3A",X"AA",X"30",
		X"DD",X"E3",X"AF",X"DD",X"ED",X"33",X"AB",X"DD",X"FE",X"DD",X"2E",X"03",X"00",X"DF",X"DD",X"D0",
		X"B0",X"00",X"DF",X"DD",X"FB",X"B0",X"0D",X"DD",X"AA",X"BB",X"D0",X"00",X"70",X"A7",X"BD",X"22",
		X"90",X"09",X"AA",X"DD",X"80",X"08",X"0A",X"24",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"00",X"00",X"22",X"00",X"00",X"0E",X"BB",X"00",X"4C",X"EC",X"00",X"2B",X"04",X"C1",X"10",X"22",
		X"24",X"CC",X"0C",X"22",X"0A",X"AA",X"AA",X"A3",X"FF",X"AA",X"FA",X"23",X"FF",X"AB",X"B0",X"32",
		X"0F",X"22",X"23",X"0D",X"ED",X"2B",X"2B",X"DD",X"EE",X"0B",X"0B",X"22",X"EE",X"0A",X"0A",X"F0",
		X"00",X"C0",X"0C",X"C0",X"B0",X"00",X"0D",X"E0",X"AB",X"E0",X"0E",X"00",X"AA",X"E0",X"00",X"00",
		X"70",X"44",X"00",X"00",X"90",X"AA",X"60",X"00",X"80",X"07",X"45",X"0C",X"00",X"08",X"A4",X"DD",
		X"00",X"00",X"0A",X"24",X"00",X"00",X"0A",X"44",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"07",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"00",X"00",X"20",X"20",X"00",X"EE",X"EB",X"02",X"00",X"EC",X"30",X"02",X"02",X"11",X"22",X"22",
		X"44",X"1A",X"22",X"22",X"42",X"AA",X"F2",X"AA",X"00",X"AA",X"3A",X"F0",X"00",X"AB",X"00",X"D0",
		X"0E",X"2E",X"EA",X"20",X"0D",X"E2",X"EA",X"AA",X"0A",X"2A",X"DA",X"AA",X"02",X"2A",X"AA",X"00",
		X"22",X"CA",X"AA",X"00",X"22",X"AA",X"AA",X"00",X"ED",X"AA",X"AA",X"00",X"D0",X"AA",X"AA",X"99",
		X"AD",X"AA",X"AA",X"99",X"7A",X"AA",X"A9",X"99",X"07",X"CA",X"99",X"99",X"09",X"DA",X"99",X"99",
		X"08",X"DD",X"99",X"99",X"00",X"AA",X"99",X"9A",X"00",X"07",X"09",X"A2",X"00",X"09",X"DD",X"A1",
		X"00",X"08",X"AA",X"22",X"00",X"00",X"0A",X"DD",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"0F",
		X"60",X"00",X"00",X"0A",X"45",X"00",X"00",X"07",X"44",X"00",X"00",X"09",X"44",X"00",X"00",X"08",
		X"AD",X"AA",X"AA",X"99",X"7A",X"AA",X"AF",X"FF",X"07",X"CA",X"FF",X"FF",X"09",X"DA",X"FF",X"FF",
		X"08",X"DD",X"FF",X"FF",X"00",X"AA",X"9F",X"FF",X"00",X"07",X"09",X"A2",X"00",X"09",X"DD",X"A1",
		X"00",X"08",X"AA",X"22",X"00",X"00",X"0A",X"DD",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"0F",
		X"60",X"00",X"00",X"0A",X"45",X"00",X"00",X"07",X"44",X"00",X"00",X"09",X"44",X"00",X"00",X"08",
		X"AD",X"AA",X"AA",X"99",X"7A",X"AA",X"AF",X"FF",X"07",X"CA",X"FF",X"FF",X"09",X"DA",X"FF",X"EF",
		X"08",X"DD",X"EF",X"FF",X"00",X"AF",X"FF",X"FF",X"00",X"FF",X"EF",X"A2",X"00",X"FF",X"FF",X"A1",
		X"00",X"FF",X"FF",X"22",X"0F",X"FF",X"FF",X"DD",X"FF",X"FF",X"F0",X"D4",X"FB",X"FF",X"00",X"0F",
		X"6F",X"FE",X"00",X"0A",X"4F",X"FF",X"00",X"07",X"44",X"F0",X"00",X"09",X"44",X"00",X"00",X"08",
		X"00",X"0E",X"2B",X"00",X"C4",X"EB",X"B2",X"00",X"44",X"B3",X"0B",X"B0",X"44",X"22",X"20",X"2B",
		X"04",X"AD",X"22",X"22",X"DB",X"AA",X"32",X"23",X"0B",X"AA",X"23",X"33",X"DD",X"3A",X"AA",X"30",
		X"DD",X"E3",X"AF",X"DD",X"ED",X"33",X"AB",X"DD",X"FE",X"DD",X"2E",X"03",X"00",X"DF",X"DD",X"D0",
		X"B0",X"00",X"DF",X"DD",X"FB",X"B0",X"0D",X"DD",X"AA",X"BB",X"D0",X"00",X"70",X"A7",X"BD",X"22",
		X"00",X"0E",X"2B",X"00",X"C4",X"EB",X"B2",X"00",X"44",X"BC",X"0B",X"B0",X"44",X"C9",X"10",X"2B",
		X"04",X"A9",X"11",X"22",X"DB",X"AC",X"91",X"23",X"0B",X"AA",X"99",X"33",X"DD",X"3A",X"AA",X"30",
		X"DD",X"E3",X"AF",X"DD",X"ED",X"33",X"AB",X"DD",X"FE",X"DD",X"2E",X"03",X"00",X"DF",X"DD",X"D0",
		X"B0",X"00",X"DF",X"DD",X"FB",X"B0",X"0D",X"DD",X"AA",X"BB",X"D0",X"00",X"70",X"A7",X"BD",X"22",
		X"00",X"B2",X"E0",X"00",X"00",X"2B",X"BE",X"4C",X"0B",X"B0",X"CB",X"44",X"B2",X"0C",X"1C",X"44",
		X"22",X"D9",X"1C",X"40",X"32",X"19",X"AA",X"BD",X"33",X"01",X"AA",X"B0",X"03",X"AA",X"A3",X"DD",
		X"DD",X"FA",X"3E",X"DD",X"DD",X"BA",X"3A",X"DE",X"30",X"22",X"DD",X"EF",X"0D",X"DD",X"FD",X"00",
		X"DD",X"FD",X"00",X"0B",X"DD",X"D0",X"0B",X"BF",X"00",X"0D",X"BB",X"AA",X"22",X"DB",X"7A",X"07",
		X"00",X"00",X"77",X"77",X"00",X"00",X"FF",X"88",X"00",X"00",X"FF",X"88",X"00",X"00",X"FF",X"88",
		X"00",X"00",X"FF",X"88",X"00",X"00",X"FF",X"88",X"00",X"00",X"FF",X"88",X"00",X"00",X"FF",X"88",
		X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"FF",X"DD",X"00",X"00",X"FF",X"DF",
		X"00",X"00",X"FF",X"DD",X"00",X"00",X"FF",X"DF",X"00",X"00",X"DF",X"DF",X"00",X"00",X"77",X"77",
		X"77",X"77",X"77",X"77",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"DF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"DF",X"DF",X"FF",X"FF",X"DF",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"88",X"88",X"8F",X"FF",X"88",X"88",X"8F",X"FF",X"88",X"88",X"8F",X"FF",
		X"88",X"88",X"8F",X"FF",X"88",X"88",X"8F",X"FF",X"88",X"88",X"8F",X"FF",X"88",X"88",X"8F",X"FF",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"DF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",
		X"DF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"DD",X"DF",X"FF",X"FF",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"FF",X"F8",X"88",X"88",X"FF",X"F8",X"88",X"88",X"FF",X"F8",X"88",X"88",
		X"FF",X"F8",X"88",X"88",X"FF",X"F8",X"88",X"88",X"FF",X"F8",X"88",X"88",X"FF",X"F8",X"88",X"88",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"DF",X"DF",X"DD",X"FF",X"DF",X"FF",X"DF",X"FF",
		X"DF",X"FF",X"DD",X"FF",X"DF",X"FF",X"DF",X"FF",X"DD",X"DF",X"DD",X"FF",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"FF",X"DD",X"DF",X"DF",X"FF",X"DF",X"DF",X"DF",
		X"FF",X"DD",X"DF",X"DF",X"FF",X"FF",X"DF",X"DF",X"FF",X"DD",X"DF",X"DD",X"77",X"77",X"77",X"77",
		X"77",X"77",X"00",X"00",X"88",X"FF",X"00",X"00",X"88",X"FF",X"00",X"00",X"88",X"FF",X"00",X"00",
		X"88",X"FF",X"00",X"00",X"88",X"FF",X"00",X"00",X"88",X"FF",X"00",X"00",X"88",X"FF",X"00",X"00",
		X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"77",X"77",X"00",X"00",
		X"44",X"00",X"00",X"44",X"45",X"00",X"00",X"54",X"67",X"00",X"00",X"76",X"09",X"00",X"00",X"90",
		X"09",X"00",X"00",X"90",X"08",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"00",X"00",X"02",X"12",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",
		X"44",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"67",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"03",X"08",X"00",X"00",X"21",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"73",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"90",X"50",X"00",X"00",X"80",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"44",X"45",X"00",X"00",X"54",X"67",X"00",X"00",X"76",X"09",X"00",X"00",X"90",
		X"09",X"00",X"60",X"90",X"08",X"05",X"45",X"80",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"60",X"05",X"44",X"44",X"45",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"45",X"75",X"44",X"44",X"67",X"07",X"44",X"44",X"09",X"09",X"44",
		X"44",X"60",X"00",X"44",X"44",X"45",X"00",X"54",X"44",X"44",X"00",X"76",X"44",X"44",X"00",X"90",
		X"44",X"44",X"60",X"90",X"75",X"44",X"45",X"80",X"07",X"44",X"44",X"00",X"09",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"05",X"44",X"45",X"00",X"44",X"44",X"67",X"00",X"44",X"44",X"09",X"00",
		X"44",X"44",X"00",X"00",X"44",X"45",X"00",X"05",X"44",X"67",X"00",X"44",X"44",X"09",X"00",X"44",
		X"44",X"60",X"00",X"44",X"44",X"45",X"05",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"75",X"44",X"44",X"45",X"07",X"44",X"44",X"69",X"09",X"44",X"44",X"09",
		X"00",X"44",X"44",X"08",X"00",X"75",X"45",X"00",X"00",X"07",X"67",X"00",X"00",X"09",X"09",X"00",
		X"00",X"00",X"09",X"00",X"50",X"00",X"08",X"05",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",
		X"44",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"67",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"60",X"00",X"08",X"05",X"45",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"60",X"05",X"44",X"44",X"45",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"45",X"75",X"44",X"44",X"67",X"07",X"44",X"44",X"09",X"09",X"44",
		X"44",X"60",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",
		X"44",X"44",X"60",X"00",X"75",X"44",X"45",X"00",X"07",X"44",X"44",X"00",X"09",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"05",X"44",X"45",X"00",X"44",X"44",X"67",X"00",X"44",X"44",X"09",X"00",
		X"44",X"44",X"00",X"00",X"44",X"45",X"00",X"05",X"44",X"67",X"00",X"44",X"44",X"09",X"00",X"44",
		X"44",X"60",X"00",X"44",X"44",X"45",X"00",X"54",X"44",X"44",X"00",X"76",X"44",X"44",X"00",X"90",
		X"44",X"44",X"60",X"90",X"75",X"44",X"45",X"80",X"07",X"44",X"44",X"00",X"09",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"05",X"44",X"45",X"00",X"44",X"44",X"67",X"00",X"44",X"44",X"09",X"00",
		X"44",X"44",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"67",X"00",X"00",X"44",X"09",X"00",X"00",
		X"44",X"60",X"00",X"44",X"44",X"45",X"05",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"75",X"44",X"44",X"45",X"07",X"44",X"44",X"69",X"09",X"44",X"44",X"09",
		X"00",X"44",X"44",X"08",X"00",X"75",X"45",X"00",X"00",X"07",X"67",X"00",X"00",X"09",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"08",X"05",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"44",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"67",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"05",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",
		X"44",X"00",X"00",X"44",X"45",X"00",X"00",X"54",X"67",X"00",X"00",X"76",X"09",X"00",X"00",X"90",
		X"09",X"00",X"00",X"90",X"08",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"44",X"45",X"00",X"00",X"54",X"67",X"00",X"00",X"76",X"09",X"00",X"00",X"90",
		X"09",X"00",X"00",X"90",X"08",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"05",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",
		X"44",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"67",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"05",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",
		X"44",X"00",X"00",X"44",X"45",X"00",X"00",X"54",X"67",X"00",X"00",X"76",X"09",X"00",X"00",X"90",
		X"09",X"00",X"00",X"90",X"08",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"44",X"45",X"00",X"05",X"44",X"67",X"00",X"44",X"44",X"09",X"00",X"44",X"44",
		X"09",X"00",X"44",X"44",X"08",X"05",X"44",X"45",X"00",X"44",X"44",X"69",X"00",X"44",X"44",X"09",
		X"00",X"44",X"44",X"68",X"05",X"44",X"44",X"45",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"45",X"75",X"44",X"44",X"67",X"07",X"44",X"44",X"09",X"09",X"44",
		X"44",X"00",X"06",X"44",X"44",X"50",X"54",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"54",X"44",X"44",X"57",X"76",X"44",X"44",X"70",X"90",X"44",X"44",X"90",
		X"90",X"44",X"44",X"00",X"80",X"54",X"44",X"50",X"00",X"76",X"44",X"44",X"00",X"90",X"44",X"44",
		X"00",X"90",X"44",X"44",X"50",X"80",X"54",X"44",X"44",X"00",X"96",X"44",X"44",X"00",X"90",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"05",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"05",X"44",X"45",X"00",X"44",X"44",X"67",X"00",X"44",X"44",X"09",
		X"00",X"44",X"44",X"09",X"05",X"44",X"45",X"08",X"44",X"44",X"69",X"00",X"44",X"44",X"09",X"00",
		X"44",X"44",X"08",X"00",X"44",X"45",X"00",X"05",X"44",X"69",X"00",X"44",X"44",X"09",X"00",X"44",
		X"44",X"00",X"00",X"44",X"45",X"00",X"05",X"44",X"67",X"00",X"44",X"44",X"09",X"00",X"44",X"44",
		X"09",X"00",X"44",X"44",X"08",X"05",X"44",X"45",X"00",X"44",X"44",X"67",X"00",X"44",X"44",X"09",
		X"00",X"44",X"44",X"09",X"05",X"44",X"45",X"08",X"44",X"44",X"69",X"00",X"44",X"44",X"09",X"00",
		X"44",X"44",X"08",X"00",X"44",X"45",X"00",X"00",X"44",X"69",X"00",X"00",X"44",X"09",X"00",X"00",
		X"44",X"00",X"00",X"44",X"45",X"00",X"05",X"44",X"67",X"00",X"44",X"44",X"09",X"00",X"44",X"44",
		X"09",X"00",X"44",X"44",X"08",X"05",X"44",X"45",X"00",X"44",X"44",X"67",X"00",X"44",X"44",X"09",
		X"00",X"44",X"44",X"09",X"05",X"44",X"45",X"08",X"44",X"44",X"69",X"00",X"44",X"44",X"09",X"00",
		X"44",X"44",X"08",X"00",X"44",X"45",X"00",X"05",X"44",X"69",X"00",X"44",X"44",X"09",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"05",X"45",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"60",X"05",X"44",X"44",X"45",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"45",X"75",X"44",X"44",X"67",X"07",X"44",X"44",X"09",X"09",X"44",
		X"44",X"60",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",
		X"44",X"44",X"60",X"00",X"75",X"44",X"45",X"00",X"07",X"44",X"44",X"00",X"09",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"05",X"44",X"45",X"00",X"44",X"44",X"67",X"00",X"44",X"44",X"09",X"00",
		X"44",X"44",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"67",X"00",X"00",X"44",X"09",X"00",X"00",
		X"44",X"60",X"00",X"44",X"44",X"45",X"05",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"75",X"44",X"44",X"45",X"07",X"44",X"44",X"69",X"09",X"44",X"44",X"09",
		X"00",X"44",X"44",X"08",X"00",X"75",X"45",X"00",X"00",X"07",X"67",X"00",X"00",X"09",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"44",X"00",X"00",X"05",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"05",X"44",X"45",X"00",X"44",X"44",X"67",X"00",X"44",X"44",X"09",
		X"00",X"44",X"44",X"09",X"05",X"44",X"45",X"08",X"44",X"44",X"69",X"00",X"44",X"44",X"09",X"00",
		X"44",X"44",X"08",X"00",X"44",X"45",X"00",X"00",X"44",X"69",X"00",X"00",X"44",X"09",X"00",X"00",
		X"44",X"60",X"00",X"44",X"44",X"45",X"05",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"75",X"44",X"44",X"45",X"07",X"44",X"44",X"67",X"09",X"44",X"44",X"00",
		X"00",X"44",X"44",X"60",X"05",X"44",X"44",X"45",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"45",X"75",X"44",X"44",X"67",X"07",X"44",X"44",X"00",X"09",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"05",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"05",X"44",X"45",X"00",X"44",X"44",X"69",X"00",X"44",X"44",X"09",
		X"00",X"44",X"44",X"68",X"05",X"44",X"44",X"45",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"45",X"75",X"44",X"44",X"67",X"07",X"44",X"44",X"09",X"09",X"44",
		X"44",X"60",X"00",X"44",X"44",X"45",X"05",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"75",X"44",X"44",X"45",X"07",X"44",X"44",X"67",X"09",X"44",X"44",X"09",
		X"00",X"44",X"44",X"09",X"05",X"44",X"45",X"08",X"44",X"44",X"67",X"00",X"44",X"44",X"09",X"00",
		X"44",X"44",X"09",X"00",X"44",X"45",X"08",X"00",X"44",X"69",X"00",X"00",X"44",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"44",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"67",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"54",X"50",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"54",X"44",X"00",X"00",X"76",X"44",X"00",X"00",X"90",X"44",
		X"00",X"00",X"FD",X"00",X"00",X"00",X"DC",X"00",X"00",X"00",X"DC",X"00",X"00",X"00",X"FC",X"00",
		X"00",X"00",X"0C",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0C",X"00",X"00",X"00",X"5C",X"50",X"00",X"00",X"0C",X"04",X"00",X"00",X"0D",X"00",
		X"00",X"00",X"0B",X"04",X"00",X"00",X"50",X"44",X"00",X"00",X"76",X"44",X"00",X"00",X"90",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"CB",X"00",X"00",X"00",X"DC",X"00",
		X"00",X"00",X"AE",X"B0",X"00",X"00",X"F0",X"A0",X"00",X"00",X"FA",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"21",X"20",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",
		X"11",X"11",X"00",X"00",X"21",X"11",X"20",X"00",X"73",X"11",X"11",X"00",X"90",X"11",X"11",X"00",
		X"0F",X"F0",X"00",X"00",X"0D",X"F0",X"00",X"00",X"0D",X"F0",X"00",X"00",X"0F",X"F0",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"24",X"20",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",
		X"10",X"00",X"00",X"00",X"21",X"11",X"20",X"00",X"73",X"11",X"11",X"00",X"90",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"00",X"D0",X"B0",X"00",X"00",X"CF",X"F0",X"00",X"00",X"EC",X"F0",X"00",X"00",
		X"DC",X"F0",X"00",X"00",X"DC",X"F0",X"00",X"00",X"BC",X"F0",X"00",X"00",X"BD",X"F0",X"00",X"00",
		X"FA",X"DB",X"00",X"00",X"FF",X"CA",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"03",X"00",X"0D",X"00",X"02",X"00",X"0D",X"D0",X"03",
		X"00",X"DD",X"D0",X"0B",X"00",X"D0",X"3D",X"05",X"00",X"00",X"2B",X"FD",X"00",X"00",X"30",X"FD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"0D",X"00",X"00",X"D0",X"0D",X"00",X"00",X"C0",X"00",X"00",X"00",X"3D",X"00",
		X"00",X"00",X"30",X"00",X"00",X"00",X"D0",X"05",X"00",X"00",X"00",X"FD",X"00",X"0D",X"D0",X"FD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"D0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0D",X"0D",X"00",X"F2",X"0C",X"0D",X"D0",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"0C",X"D0",X"FD",X"00",X"03",X"30",X"FD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"03",
		X"00",X"0D",X"30",X"03",X"00",X"03",X"20",X"0D",X"00",X"D2",X"2D",X"FD",X"00",X"0D",X"D2",X"FD",
		X"00",X"D0",X"00",X"DC",X"00",X"D0",X"D5",X"DF",X"0D",X"3D",X"DF",X"FF",X"D2",X"23",X"DD",X"FF",
		X"D2",X"22",X"BD",X"FF",X"DB",X"D3",X"3D",X"F5",X"DD",X"DD",X"FF",X"69",X"0D",X"DD",X"FF",X"09",
		X"0D",X"CC",X"FF",X"68",X"0C",X"2D",X"F4",X"45",X"DD",X"FF",X"44",X"44",X"DC",X"FF",X"44",X"44",
		X"D3",X"FF",X"44",X"44",X"DF",X"F5",X"75",X"44",X"FF",X"67",X"07",X"44",X"FF",X"09",X"09",X"44",
		X"0C",X"D3",X"D0",X"F2",X"0C",X"2D",X"C5",X"DF",X"00",X"23",X"CD",X"FF",X"00",X"C3",X"3D",X"FF",
		X"0D",X"DC",X"23",X"FF",X"0D",X"DD",X"2D",X"F5",X"0C",X"DD",X"FF",X"69",X"0D",X"DD",X"FF",X"09",
		X"0D",X"C3",X"FF",X"68",X"0D",X"2B",X"F4",X"45",X"D3",X"FF",X"44",X"44",X"D2",X"FF",X"44",X"44",
		X"D3",X"FF",X"44",X"44",X"FF",X"F5",X"75",X"44",X"FF",X"67",X"07",X"44",X"FF",X"09",X"09",X"44",
		X"00",X"DC",X"D0",X"DC",X"00",X"3D",X"3D",X"DF",X"0D",X"2D",X"2D",X"FF",X"D0",X"2D",X"23",X"FF",
		X"D0",X"BD",X"D2",X"FF",X"D0",X"3D",X"DD",X"F5",X"CD",X"C3",X"FF",X"69",X"03",X"32",X"FF",X"09",
		X"0D",X"2C",X"FF",X"68",X"0D",X"3D",X"F4",X"45",X"D3",X"FF",X"44",X"44",X"D2",X"FF",X"44",X"44",
		X"D3",X"FF",X"44",X"44",X"FF",X"F5",X"75",X"44",X"FF",X"67",X"07",X"44",X"FF",X"09",X"09",X"44",
		X"00",X"D2",X"2D",X"DD",X"00",X"B2",X"23",X"DF",X"00",X"D3",X"D2",X"FF",X"0D",X"03",X"D3",X"FF",
		X"0B",X"DB",X"DD",X"FF",X"03",X"B2",X"DD",X"F5",X"0B",X"2D",X"FF",X"69",X"0D",X"3D",X"FF",X"09",
		X"03",X"DD",X"FF",X"68",X"02",X"D3",X"F4",X"45",X"D3",X"FF",X"44",X"44",X"D3",X"FF",X"44",X"44",
		X"DC",X"FF",X"44",X"44",X"FF",X"F5",X"75",X"44",X"FF",X"67",X"07",X"44",X"FF",X"09",X"09",X"44",
		X"00",X"00",X"D3",X"DD",X"00",X"00",X"DD",X"DF",X"00",X"0D",X"DF",X"FF",X"00",X"03",X"DD",X"FF",
		X"00",X"D2",X"DD",X"FF",X"00",X"22",X"BD",X"F5",X"0C",X"33",X"FF",X"69",X"0C",X"BD",X"FF",X"09",
		X"03",X"DD",X"FF",X"68",X"0B",X"D3",X"F4",X"45",X"DC",X"FF",X"44",X"44",X"DD",X"FF",X"44",X"44",
		X"DC",X"FF",X"44",X"44",X"FF",X"F5",X"75",X"44",X"FF",X"67",X"07",X"44",X"FF",X"09",X"09",X"44",
		X"00",X"D0",X"00",X"DC",X"00",X"D0",X"D5",X"DF",X"0D",X"3D",X"DF",X"FF",X"D2",X"23",X"DD",X"FF",
		X"D2",X"22",X"BD",X"FF",X"DB",X"D3",X"3D",X"F5",X"DD",X"DD",X"FF",X"69",X"0D",X"DD",X"FF",X"09",
		X"0D",X"CC",X"FF",X"68",X"0C",X"2D",X"FF",X"F5",X"DD",X"FF",X"FF",X"FF",X"DC",X"FF",X"FF",X"FF",
		X"D3",X"FF",X"FF",X"FF",X"DF",X"F5",X"75",X"FF",X"FF",X"67",X"07",X"FF",X"FF",X"09",X"09",X"FF",
		X"0C",X"D3",X"D0",X"F2",X"0C",X"2D",X"C5",X"DF",X"00",X"23",X"CD",X"FF",X"00",X"C3",X"3D",X"FF",
		X"0D",X"DC",X"23",X"FF",X"0D",X"DD",X"2D",X"F5",X"0C",X"DD",X"FF",X"69",X"0D",X"DD",X"FF",X"09",
		X"0D",X"C3",X"FF",X"68",X"0D",X"2B",X"FF",X"F5",X"D3",X"FF",X"FF",X"FF",X"D2",X"FF",X"FF",X"FF",
		X"D3",X"FF",X"FF",X"FF",X"FF",X"F5",X"75",X"FF",X"FF",X"67",X"07",X"FF",X"FF",X"09",X"09",X"FF",
		X"00",X"DC",X"D0",X"DC",X"00",X"3D",X"3D",X"DF",X"0D",X"2D",X"2D",X"FF",X"D0",X"2D",X"23",X"FF",
		X"D0",X"BD",X"D2",X"FF",X"D0",X"3D",X"DD",X"F5",X"CD",X"C3",X"FF",X"69",X"03",X"32",X"FF",X"09",
		X"0D",X"2C",X"FF",X"68",X"0D",X"3D",X"FF",X"F5",X"D3",X"FF",X"FF",X"FF",X"D2",X"FF",X"FF",X"FF",
		X"D3",X"FF",X"FF",X"FF",X"FF",X"F5",X"75",X"FF",X"FF",X"67",X"07",X"FF",X"FF",X"09",X"09",X"FF",
		X"00",X"D2",X"2D",X"DD",X"00",X"B2",X"23",X"DF",X"00",X"D3",X"D2",X"FF",X"0D",X"03",X"D3",X"FF",
		X"0B",X"DB",X"DD",X"FF",X"03",X"B2",X"DD",X"F5",X"0B",X"2D",X"FF",X"69",X"0D",X"3D",X"FF",X"09",
		X"03",X"DD",X"FF",X"68",X"02",X"D3",X"FF",X"F5",X"D3",X"FF",X"FF",X"FF",X"D3",X"FF",X"FF",X"FF",
		X"DC",X"FF",X"FF",X"FF",X"FF",X"F5",X"75",X"FF",X"FF",X"67",X"07",X"FF",X"FF",X"09",X"09",X"FF",
		X"00",X"00",X"D3",X"DD",X"00",X"00",X"DD",X"DF",X"00",X"0D",X"DF",X"FF",X"00",X"03",X"DD",X"FF",
		X"00",X"D2",X"DD",X"FF",X"00",X"22",X"BD",X"F5",X"0C",X"33",X"FF",X"69",X"0C",X"BD",X"FF",X"09",
		X"03",X"DD",X"FF",X"68",X"0B",X"D3",X"FF",X"F5",X"DC",X"FF",X"FF",X"FF",X"DD",X"FF",X"FF",X"FF",
		X"DC",X"FF",X"FF",X"FF",X"FF",X"F5",X"75",X"FF",X"FF",X"67",X"07",X"FF",X"FF",X"09",X"09",X"FF",
		X"00",X"D0",X"00",X"DC",X"00",X"D0",X"D5",X"DF",X"0D",X"3D",X"DF",X"FF",X"D2",X"23",X"DD",X"FF",
		X"D2",X"22",X"BD",X"FF",X"DB",X"D3",X"3D",X"F5",X"DD",X"DD",X"FF",X"69",X"0D",X"DD",X"FF",X"09",
		X"0D",X"CC",X"FF",X"6D",X"0C",X"2D",X"FF",X"F3",X"DD",X"FD",X"FF",X"F2",X"DC",X"FD",X"DF",X"F3",
		X"D3",X"DD",X"DF",X"FB",X"DF",X"D5",X"3D",X"FF",X"FF",X"67",X"2B",X"FD",X"FF",X"09",X"39",X"FD",
		X"0C",X"D3",X"D0",X"F2",X"0C",X"2D",X"C5",X"DF",X"00",X"23",X"CD",X"FF",X"00",X"C3",X"3D",X"FF",
		X"0D",X"DC",X"23",X"FF",X"0D",X"DD",X"2D",X"FD",X"0C",X"DD",X"FF",X"6C",X"0D",X"DD",X"FF",X"0B",
		X"0D",X"C3",X"FF",X"6D",X"0D",X"2B",X"DF",X"FD",X"D3",X"FF",X"CF",X"FF",X"D2",X"FF",X"3D",X"FF",
		X"D3",X"FF",X"3F",X"FF",X"FF",X"F5",X"D5",X"FF",X"FF",X"67",X"07",X"FD",X"FF",X"0D",X"D9",X"FD",
		X"00",X"DC",X"D0",X"DC",X"00",X"3D",X"3D",X"DF",X"0D",X"2D",X"2D",X"FF",X"D0",X"2D",X"23",X"FD",
		X"D0",X"BD",X"D2",X"FD",X"D0",X"3D",X"DD",X"FD",X"CD",X"C3",X"FF",X"6D",X"03",X"32",X"DF",X"09",
		X"0D",X"2C",X"DF",X"68",X"0D",X"3D",X"BF",X"F5",X"D3",X"FF",X"DF",X"FF",X"D2",X"FF",X"FF",X"FF",
		X"D3",X"FF",X"FF",X"FF",X"FF",X"F5",X"75",X"FD",X"FD",X"6D",X"07",X"F2",X"FC",X"0D",X"D9",X"F3",
		X"00",X"D2",X"2D",X"DD",X"00",X"B2",X"23",X"DF",X"00",X"D3",X"D2",X"FF",X"0D",X"03",X"D3",X"FD",
		X"0B",X"DB",X"DD",X"FF",X"03",X"B2",X"DD",X"F5",X"0B",X"2D",X"DF",X"69",X"0D",X"3D",X"CF",X"09",
		X"03",X"DD",X"DF",X"68",X"02",X"D3",X"FF",X"F5",X"D3",X"FF",X"FF",X"FD",X"D3",X"FF",X"FF",X"F2",
		X"DC",X"FF",X"FF",X"F3",X"FF",X"F5",X"75",X"F3",X"FF",X"6C",X"D7",X"FD",X"FF",X"03",X"39",X"FD",
		X"00",X"00",X"D3",X"DD",X"00",X"00",X"DD",X"DF",X"00",X"0D",X"DF",X"FF",X"00",X"03",X"DD",X"FF",
		X"00",X"D2",X"DD",X"FF",X"00",X"22",X"BD",X"F5",X"0C",X"33",X"DF",X"69",X"0C",X"BD",X"FF",X"09",
		X"03",X"DD",X"FF",X"68",X"0B",X"D3",X"FF",X"FD",X"DC",X"FF",X"FF",X"F2",X"DD",X"FF",X"FF",X"F3",
		X"DC",X"FD",X"3F",X"F3",X"FF",X"F3",X"25",X"FD",X"FF",X"D2",X"2D",X"FD",X"FF",X"0D",X"D2",X"FD",
		X"FF",X"D0",X"00",X"DC",X"FF",X"D5",X"D5",X"DF",X"FD",X"3D",X"DF",X"FF",X"D2",X"23",X"DD",X"FF",
		X"D2",X"22",X"BD",X"FF",X"DB",X"D3",X"3D",X"F5",X"DD",X"DD",X"FF",X"67",X"0D",X"DD",X"FF",X"00",
		X"0D",X"CC",X"FF",X"60",X"0C",X"2D",X"F4",X"45",X"DD",X"FF",X"44",X"44",X"DC",X"FF",X"44",X"44",
		X"D3",X"FF",X"44",X"44",X"DF",X"F5",X"75",X"44",X"FF",X"67",X"07",X"44",X"FF",X"00",X"09",X"44",
		X"FC",X"D3",X"D0",X"F2",X"FC",X"2D",X"C5",X"DF",X"FF",X"23",X"CD",X"FF",X"FF",X"C3",X"3D",X"FF",
		X"FD",X"DC",X"23",X"FF",X"7D",X"DD",X"2D",X"F5",X"0C",X"DD",X"FF",X"67",X"0D",X"DD",X"FF",X"00",
		X"0D",X"C3",X"FF",X"60",X"0D",X"2B",X"F4",X"45",X"D3",X"FF",X"44",X"44",X"D2",X"FF",X"44",X"44",
		X"D3",X"FF",X"44",X"44",X"FF",X"F5",X"75",X"44",X"FF",X"67",X"07",X"44",X"FF",X"00",X"09",X"44",
		X"FF",X"DC",X"D0",X"DC",X"FF",X"3D",X"3D",X"DF",X"FD",X"2D",X"2D",X"FF",X"DF",X"2D",X"23",X"FF",
		X"DF",X"BD",X"D2",X"FF",X"D5",X"3D",X"DD",X"F5",X"CD",X"C3",X"FF",X"67",X"03",X"32",X"FF",X"00",
		X"0D",X"2C",X"FF",X"60",X"0D",X"3D",X"F4",X"45",X"D3",X"FF",X"44",X"44",X"D2",X"FF",X"44",X"44",
		X"D3",X"FF",X"44",X"44",X"FF",X"F5",X"75",X"44",X"FF",X"67",X"07",X"44",X"FF",X"00",X"09",X"44",
		X"FF",X"D2",X"2D",X"DD",X"FF",X"B2",X"23",X"DF",X"FF",X"D3",X"D2",X"FF",X"FD",X"F3",X"D3",X"FF",
		X"FB",X"DB",X"DD",X"FF",X"73",X"B2",X"DD",X"F5",X"0B",X"2D",X"FF",X"67",X"0D",X"3D",X"FF",X"00",
		X"03",X"DD",X"FF",X"60",X"02",X"D3",X"F4",X"45",X"D3",X"FF",X"44",X"44",X"D3",X"FF",X"44",X"44",
		X"DC",X"FF",X"44",X"44",X"FF",X"F5",X"75",X"44",X"FF",X"67",X"07",X"44",X"FF",X"00",X"09",X"44",
		X"FF",X"60",X"D3",X"DD",X"FF",X"F5",X"DD",X"DF",X"FF",X"FD",X"DF",X"FF",X"FF",X"F3",X"DD",X"FF",
		X"FF",X"D2",X"DD",X"FF",X"75",X"22",X"BD",X"F5",X"0C",X"33",X"FF",X"67",X"0C",X"BD",X"FF",X"00",
		X"03",X"DD",X"FF",X"60",X"0B",X"D3",X"F4",X"45",X"DC",X"FF",X"44",X"44",X"DD",X"FF",X"44",X"44",
		X"DC",X"FF",X"44",X"44",X"FF",X"F5",X"75",X"44",X"FF",X"67",X"07",X"44",X"FF",X"00",X"09",X"44",
		X"FF",X"D0",X"00",X"DC",X"FF",X"D5",X"D5",X"DF",X"FD",X"3D",X"DF",X"FF",X"D2",X"23",X"DD",X"FF",
		X"D2",X"22",X"BD",X"FF",X"DB",X"D3",X"3D",X"F5",X"DD",X"DD",X"FF",X"67",X"0D",X"DD",X"FF",X"00",
		X"0D",X"CC",X"FF",X"60",X"0C",X"2D",X"FF",X"F5",X"DD",X"FF",X"FF",X"FF",X"DC",X"FF",X"FF",X"FF",
		X"D3",X"FF",X"FF",X"FF",X"DF",X"F5",X"75",X"FF",X"FF",X"67",X"07",X"FF",X"FF",X"00",X"09",X"FF",
		X"FC",X"D3",X"D0",X"F2",X"FC",X"2D",X"C5",X"DF",X"FF",X"23",X"CD",X"FF",X"FF",X"C3",X"3D",X"FF",
		X"FD",X"DC",X"23",X"FF",X"7D",X"DD",X"2D",X"F5",X"0C",X"DD",X"FF",X"67",X"0D",X"DD",X"FF",X"00",
		X"0D",X"C3",X"FF",X"60",X"0D",X"2B",X"FF",X"F5",X"D3",X"FF",X"FF",X"FF",X"D2",X"FF",X"FF",X"FF",
		X"D3",X"FF",X"FF",X"FF",X"FF",X"F5",X"75",X"FF",X"FF",X"67",X"07",X"FF",X"FF",X"00",X"09",X"FF",
		X"FF",X"DC",X"D0",X"DC",X"FF",X"3D",X"3D",X"DF",X"FD",X"2D",X"2D",X"FF",X"DF",X"2D",X"23",X"FF",
		X"DF",X"BD",X"D2",X"FF",X"D5",X"3D",X"DD",X"F5",X"CD",X"C3",X"FF",X"67",X"03",X"32",X"FF",X"00",
		X"0D",X"2C",X"FF",X"60",X"0D",X"3D",X"FF",X"F5",X"D3",X"FF",X"FF",X"FF",X"D2",X"FF",X"FF",X"FF",
		X"D3",X"FF",X"FF",X"FF",X"FF",X"F5",X"75",X"FF",X"FF",X"67",X"07",X"FF",X"FF",X"00",X"09",X"FF",
		X"FF",X"D2",X"2D",X"DD",X"FF",X"B2",X"23",X"DF",X"FF",X"D3",X"D2",X"FF",X"FD",X"F3",X"D3",X"FF",
		X"FB",X"DB",X"DD",X"FF",X"73",X"B2",X"DD",X"F5",X"0B",X"2D",X"FF",X"67",X"0D",X"3D",X"FF",X"00",
		X"03",X"DD",X"FF",X"60",X"02",X"D3",X"FF",X"F5",X"D3",X"FF",X"FF",X"FF",X"D3",X"FF",X"FF",X"FF",
		X"DC",X"FF",X"FF",X"FF",X"FF",X"F5",X"75",X"FF",X"FF",X"67",X"07",X"FF",X"FF",X"00",X"09",X"FF",
		X"FF",X"60",X"D3",X"DD",X"FF",X"F5",X"DD",X"DF",X"FF",X"FD",X"DF",X"FF",X"FF",X"F3",X"DD",X"FF",
		X"FF",X"D2",X"DD",X"FF",X"75",X"22",X"BD",X"F5",X"0C",X"33",X"FF",X"67",X"0C",X"BD",X"FF",X"00",
		X"03",X"DD",X"FF",X"60",X"0B",X"D3",X"FF",X"F5",X"DC",X"FF",X"FF",X"FF",X"DD",X"FF",X"FF",X"FF",
		X"DC",X"FF",X"FF",X"FF",X"FF",X"F5",X"75",X"FF",X"FF",X"67",X"07",X"FF",X"FF",X"00",X"09",X"FF",
		X"FF",X"D0",X"00",X"DC",X"FF",X"D5",X"D5",X"DF",X"FD",X"3D",X"DF",X"FF",X"D2",X"23",X"DD",X"FF",
		X"D2",X"22",X"BD",X"FF",X"DB",X"D3",X"3D",X"F5",X"DD",X"DD",X"FF",X"67",X"0D",X"DD",X"FF",X"00",
		X"0D",X"CC",X"FF",X"6D",X"0C",X"2D",X"FF",X"F3",X"DD",X"FD",X"FF",X"F2",X"DC",X"FD",X"DF",X"F3",
		X"D3",X"DD",X"DF",X"FB",X"DF",X"D5",X"3D",X"FF",X"FF",X"67",X"2B",X"FD",X"FF",X"00",X"39",X"FD",
		X"FC",X"D3",X"D0",X"F2",X"FC",X"2D",X"C5",X"DF",X"FF",X"23",X"CD",X"FF",X"FF",X"C3",X"3D",X"FF",
		X"FD",X"DC",X"23",X"FF",X"7D",X"DD",X"2D",X"FD",X"0C",X"DD",X"FF",X"6C",X"0D",X"DD",X"FF",X"0B",
		X"0D",X"C3",X"FF",X"6D",X"0D",X"2B",X"DF",X"FD",X"D3",X"FF",X"CF",X"FF",X"D2",X"FF",X"3D",X"FF",
		X"D3",X"FF",X"3F",X"FF",X"FF",X"F5",X"D5",X"FF",X"FF",X"67",X"07",X"FD",X"FF",X"0D",X"D9",X"FD",
		X"FF",X"DC",X"D0",X"DC",X"FF",X"3D",X"3D",X"DF",X"FD",X"2D",X"2D",X"FF",X"DF",X"2D",X"23",X"FD",
		X"DF",X"BD",X"D2",X"FD",X"D5",X"3D",X"DD",X"FD",X"CD",X"C3",X"FF",X"6D",X"03",X"32",X"DF",X"00",
		X"0D",X"2C",X"DF",X"60",X"0D",X"3D",X"BF",X"F5",X"D3",X"FF",X"DF",X"FF",X"D2",X"FF",X"FF",X"FF",
		X"D3",X"FF",X"FF",X"FF",X"FF",X"F5",X"75",X"FD",X"FD",X"6D",X"07",X"F2",X"FC",X"0D",X"D9",X"F3",
		X"FF",X"D2",X"2D",X"DD",X"FF",X"B2",X"23",X"DF",X"FF",X"D3",X"D2",X"FF",X"FD",X"F3",X"D3",X"FD",
		X"FB",X"DB",X"DD",X"FF",X"73",X"B2",X"DD",X"F5",X"0B",X"2D",X"DF",X"67",X"0D",X"3D",X"CF",X"00",
		X"03",X"DD",X"DF",X"60",X"02",X"D3",X"FF",X"F5",X"D3",X"FF",X"FF",X"FD",X"D3",X"FF",X"FF",X"F2",
		X"DC",X"FF",X"FF",X"F3",X"FF",X"F5",X"75",X"F3",X"FF",X"6C",X"D7",X"FD",X"FF",X"03",X"39",X"FD",
		X"FF",X"60",X"D3",X"DD",X"FF",X"F5",X"DD",X"DF",X"FF",X"FD",X"DF",X"FF",X"FF",X"F3",X"DD",X"FF",
		X"FF",X"D2",X"DD",X"FF",X"75",X"22",X"BD",X"F5",X"0C",X"33",X"DF",X"67",X"0C",X"BD",X"FF",X"00",
		X"03",X"DD",X"FF",X"60",X"0B",X"D3",X"FF",X"FD",X"DC",X"FF",X"FF",X"F2",X"DD",X"FF",X"FF",X"F3",
		X"DC",X"FD",X"3F",X"F3",X"FF",X"F3",X"25",X"FD",X"FF",X"D2",X"2D",X"FD",X"FF",X"0D",X"D2",X"FD",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"05",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"05",X"FF",X"F5",X"00",X"FF",X"FF",X"69",X"00",X"FF",X"FF",X"09",
		X"00",X"FF",X"FF",X"68",X"05",X"FF",X"F4",X"45",X"FF",X"FF",X"44",X"44",X"FF",X"FF",X"44",X"44",
		X"FF",X"FF",X"44",X"44",X"FF",X"F5",X"75",X"44",X"FF",X"67",X"07",X"44",X"FF",X"09",X"09",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"FF",X"60",X"00",X"44",X"FF",X"45",X"05",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"75",X"44",X"44",X"45",X"07",X"44",X"44",X"67",X"09",X"44",X"44",X"00",
		X"00",X"44",X"44",X"60",X"05",X"44",X"44",X"45",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"45",X"75",X"44",X"44",X"67",X"07",X"44",X"44",X"00",X"09",X"44",
		X"FF",X"60",X"00",X"FF",X"FF",X"F5",X"05",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"75",X"FF",X"FF",X"F5",X"07",X"FF",X"FF",X"67",X"09",X"FF",X"FF",X"00",
		X"00",X"FF",X"FF",X"60",X"05",X"FF",X"F4",X"45",X"FF",X"FF",X"44",X"44",X"FF",X"FF",X"44",X"44",
		X"FF",X"FF",X"44",X"44",X"FF",X"F5",X"75",X"44",X"FF",X"67",X"07",X"44",X"FF",X"00",X"09",X"44",
		X"FF",X"60",X"00",X"FF",X"FF",X"F5",X"05",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"75",X"FF",X"FF",X"F5",X"07",X"FF",X"FF",X"67",X"09",X"FF",X"FF",X"00",
		X"00",X"FF",X"FF",X"60",X"05",X"FF",X"FF",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"75",X"FF",X"FF",X"67",X"07",X"FF",X"FF",X"00",X"09",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
