library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity inferno_graph3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of inferno_graph3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"31",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"31",X"11",X"13",X"00",X"11",X"11",X"77",X"00",X"11",X"11",X"09",X"00",X"11",X"11",X"00",
		X"31",X"11",X"13",X"00",X"11",X"11",X"77",X"00",X"11",X"11",X"09",X"00",X"11",X"11",X"00",X"00",
		X"11",X"13",X"00",X"00",X"11",X"77",X"00",X"00",X"11",X"09",X"00",X"00",X"11",X"00",X"00",X"00",
		X"13",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"13",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"13",X"00",X"00",X"11",X"77",X"00",X"00",X"31",X"09",X"00",X"00",X"07",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"11",X"13",X"00",X"00",X"11",X"11",X"00",X"00",X"11",
		X"11",X"00",X"31",X"11",X"11",X"00",X"11",X"11",X"11",X"13",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"13",X"11",X"11",X"11",X"77",X"31",X"11",X"11",X"09",X"07",X"11",X"11",X"00",
		X"31",X"11",X"13",X"00",X"11",X"11",X"77",X"00",X"11",X"11",X"09",X"00",X"11",X"11",X"00",X"00",
		X"11",X"13",X"00",X"00",X"11",X"77",X"00",X"00",X"11",X"09",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"13",X"00",X"00",X"11",X"11",X"00",X"00",
		X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"31",X"11",X"13",X"00",X"07",X"11",X"11",X"00",
		X"31",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"13",X"11",X"11",X"11",X"11",
		X"11",X"13",X"11",X"11",X"11",X"77",X"11",X"11",X"11",X"00",X"31",X"11",X"11",X"00",X"07",X"11",
		X"13",X"00",X"09",X"11",X"77",X"00",X"00",X"11",X"09",X"00",X"00",X"31",X"00",X"00",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"31",X"11",X"13",X"00",X"11",X"11",X"77",X"00",X"11",X"11",X"09",X"00",X"11",X"11",X"00",X"00",
		X"11",X"13",X"00",X"31",X"11",X"77",X"00",X"11",X"11",X"09",X"00",X"11",X"11",X"00",X"00",X"11",
		X"13",X"00",X"31",X"11",X"77",X"00",X"11",X"11",X"09",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"31",X"11",X"13",X"00",X"11",X"11",X"77",X"00",X"11",X"11",X"09",X"00",X"11",X"11",X"00",
		X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"31",X"11",X"13",X"00",X"07",X"11",X"11",
		X"00",X"09",X"11",X"11",X"00",X"00",X"11",X"11",X"13",X"00",X"31",X"11",X"11",X"00",X"07",X"11",
		X"11",X"00",X"31",X"11",X"11",X"00",X"11",X"11",X"11",X"13",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"13",X"11",X"11",X"11",X"77",X"31",X"11",X"11",X"00",X"07",X"11",X"11",X"00",
		X"31",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"13",X"11",X"11",X"11",X"11",
		X"11",X"13",X"11",X"11",X"11",X"77",X"11",X"11",X"11",X"90",X"31",X"11",X"11",X"90",X"07",X"11",
		X"11",X"80",X"09",X"11",X"11",X"00",X"00",X"11",X"11",X"13",X"00",X"31",X"11",X"11",X"00",X"07",
		X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"31",X"11",X"13",X"00",X"07",X"11",X"11",X"00",
		X"31",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"13",X"11",X"11",X"11",X"11",
		X"11",X"13",X"11",X"11",X"11",X"77",X"11",X"11",X"11",X"90",X"31",X"11",X"11",X"90",X"07",X"11",
		X"11",X"80",X"31",X"11",X"11",X"00",X"11",X"11",X"11",X"13",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"13",X"11",X"11",X"11",X"77",X"31",X"11",X"11",X"00",X"07",X"11",X"11",X"00",
		X"00",X"11",X"13",X"00",X"00",X"11",X"77",X"00",X"00",X"31",X"09",X"00",X"00",X"07",X"00",X"00",
		X"00",X"09",X"00",X"31",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"31",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"31",X"11",X"13",X"00",X"11",X"11",X"77",X"00",X"11",X"11",X"09",X"00",X"11",X"11",X"00",
		X"07",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"30",X"00",X"72",X"11",X"12",
		X"00",X"97",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"72",X"11",
		X"00",X"00",X"07",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"72",
		X"00",X"31",X"00",X"07",X"00",X"11",X"00",X"00",X"00",X"11",X"13",X"00",X"00",X"11",X"11",X"00",
		X"00",X"11",X"13",X"00",X"00",X"11",X"77",X"00",X"00",X"31",X"09",X"00",X"00",X"07",X"00",X"02",
		X"00",X"09",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"02",X"11",
		X"00",X"00",X"07",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"72",
		X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"13",X"00",X"00",X"11",X"77",X"00",X"00",X"31",X"09",X"00",X"00",X"07",X"00",X"00",
		X"00",X"09",X"00",X"31",X"00",X"00",X"00",X"11",X"13",X"00",X"00",X"11",X"11",X"00",X"00",X"11",
		X"11",X"00",X"31",X"11",X"11",X"00",X"11",X"11",X"11",X"13",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"13",X"11",X"11",X"11",X"77",X"31",X"11",X"11",X"09",X"07",X"11",X"11",X"00",
		X"07",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"30",X"00",X"72",X"11",X"12",
		X"00",X"97",X"11",X"11",X"00",X"00",X"11",X"11",X"13",X"00",X"11",X"11",X"11",X"00",X"72",X"11",
		X"13",X"00",X"11",X"11",X"77",X"00",X"11",X"11",X"09",X"00",X"11",X"11",X"00",X"02",X"11",X"12",
		X"00",X"11",X"11",X"37",X"00",X"11",X"11",X"90",X"00",X"11",X"11",X"90",X"02",X"11",X"12",X"80",
		X"31",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"13",X"11",X"11",X"11",X"11",
		X"11",X"13",X"11",X"11",X"11",X"77",X"11",X"11",X"11",X"00",X"31",X"11",X"11",X"00",X"07",X"11",
		X"13",X"00",X"09",X"11",X"77",X"00",X"00",X"11",X"09",X"00",X"00",X"31",X"00",X"00",X"00",X"07",
		X"00",X"31",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"13",X"00",X"00",X"11",X"11",X"00",
		X"46",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"31",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"31",X"11",X"13",X"00",X"11",X"11",X"77",X"00",X"11",X"11",X"09",X"00",X"11",X"11",X"00",
		X"07",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"30",X"00",X"72",X"11",X"12",
		X"00",X"97",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"72",X"11",
		X"00",X"00",X"07",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"72",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"45",X"00",X"00",X"00",
		X"46",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"02",X"11",
		X"00",X"00",X"07",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"72",
		X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"46",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",
		X"31",X"00",X"00",X"31",X"11",X"00",X"00",X"11",X"13",X"00",X"00",X"11",X"77",X"11",X"00",X"11",
		X"77",X"13",X"31",X"11",X"77",X"77",X"11",X"11",X"31",X"77",X"11",X"11",X"11",X"77",X"11",X"11",
		X"99",X"31",X"11",X"13",X"00",X"11",X"11",X"97",X"00",X"11",X"11",X"90",X"00",X"11",X"11",X"80",
		X"31",X"11",X"13",X"00",X"11",X"11",X"77",X"00",X"11",X"11",X"77",X"00",X"11",X"11",X"77",X"00",
		X"11",X"13",X"64",X"00",X"11",X"77",X"44",X"00",X"11",X"00",X"46",X"00",X"11",X"00",X"77",X"44",
		X"13",X"00",X"77",X"46",X"77",X"00",X"77",X"77",X"09",X"00",X"64",X"77",X"00",X"00",X"44",X"77",
		X"00",X"00",X"99",X"64",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"46",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",
		X"31",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"13",X"00",X"00",X"00",X"77",X"11",X"00",X"00",
		X"77",X"13",X"00",X"00",X"77",X"77",X"00",X"00",X"31",X"77",X"00",X"00",X"11",X"77",X"00",X"00",
		X"99",X"31",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"13",X"00",X"00",X"11",X"11",X"00",
		X"00",X"11",X"13",X"00",X"00",X"11",X"77",X"00",X"00",X"31",X"77",X"00",X"00",X"09",X"77",X"00",
		X"00",X"09",X"64",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"46",X"00",X"00",X"00",X"77",X"44",
		X"00",X"00",X"77",X"46",X"00",X"00",X"77",X"77",X"00",X"00",X"64",X"77",X"00",X"00",X"44",X"77",
		X"00",X"00",X"99",X"64",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"02",X"22",X"00",X"01",X"44",X"0B",X"2B",X"02",X"24",X"CC",X"22",X"0E",X"40",X"11",X"B2",X"B3",
		X"0A",X"11",X"0B",X"B3",X"F2",X"11",X"00",X"3E",X"FF",X"AC",X"C1",X"EE",X"BB",X"AA",X"A0",X"EE",
		X"DD",X"AA",X"AB",X"EF",X"DD",X"33",X"F2",X"DD",X"DD",X"AA",X"E2",X"DD",X"CE",X"DD",X"BB",X"DD",
		X"D0",X"DD",X"DD",X"DD",X"BB",X"00",X"DD",X"20",X"0A",X"BB",X"01",X"00",X"0A",X"0A",X"D2",X"D0",
		X"00",X"00",X"4D",X"DD",X"00",X"00",X"7A",X"4D",X"00",X"00",X"90",X"42",X"00",X"00",X"80",X"A4",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"46",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"00",X"EE",X"B0",X"00",X"02",X"EB",X"22",X"01",X"D4",X"CC",X"B2",X"0E",X"40",X"11",X"0B",X"B3",
		X"0A",X"11",X"10",X"BE",X"3A",X"AA",X"A0",X"3E",X"33",X"AA",X"BB",X"EE",X"33",X"AA",X"22",X"EF",
		X"FE",X"BB",X"22",X"DD",X"DD",X"22",X"F3",X"DD",X"DD",X"22",X"22",X"DA",X"F0",X"FF",X"BF",X"F0",
		X"00",X"0C",X"0C",X"C0",X"E0",X"0C",X"00",X"00",X"B0",X"0E",X"00",X"00",X"0A",X"20",X"20",X"00",
		X"0A",X"D0",X"C0",X"00",X"0A",X"44",X"10",X"D0",X"00",X"0A",X"DD",X"20",X"00",X"00",X"4D",X"DD",
		X"00",X"00",X"A4",X"4D",X"00",X"00",X"7A",X"42",X"00",X"00",X"90",X"A4",X"00",X"00",X"80",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"46",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EB",X"22",X"B0",X"00",X"1C",X"22",X"ED",X"44",X"00",X"AB",X"2D",
		X"40",X"0A",X"22",X"23",X"00",X"A2",X"2A",X"A0",X"0A",X"22",X"FF",X"F0",X"EA",X"22",X"FC",X"C0",
		X"3A",X"F3",X"AD",X"AA",X"3A",X"20",X"AA",X"AA",X"32",X"CC",X"AA",X"AA",X"22",X"AC",X"AA",X"AA",
		X"22",X"A2",X"A0",X"0A",X"2A",X"AA",X"A0",X"0A",X"DA",X"AA",X"A0",X"07",X"0A",X"AA",X"AA",X"00",
		X"D0",X"AA",X"99",X"90",X"AD",X"AA",X"99",X"9A",X"0A",X"AD",X"99",X"9A",X"0A",X"A2",X"D9",X"9A",
		X"0A",X"0C",X"C9",X"AA",X"00",X"DD",X"19",X"9A",X"00",X"0A",X"19",X"AA",X"00",X"0A",X"2C",X"AA",
		X"00",X"00",X"DD",X"D0",X"00",X"00",X"A7",X"DD",X"00",X"00",X"7A",X"4D",X"00",X"00",X"90",X"42",
		X"00",X"00",X"80",X"A4",X"00",X"00",X"00",X"A0",X"46",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"D0",X"AA",X"9F",X"90",X"AD",X"AA",X"FF",X"9A",X"0A",X"AD",X"FF",X"FA",X"0A",X"A2",X"FF",X"FF",
		X"0A",X"0C",X"FF",X"FA",X"00",X"DD",X"FF",X"9A",X"00",X"0A",X"FF",X"AA",X"00",X"0A",X"2C",X"AA",
		X"00",X"00",X"DD",X"D0",X"00",X"00",X"A7",X"DD",X"00",X"00",X"7A",X"4D",X"00",X"00",X"90",X"42",
		X"00",X"00",X"80",X"A4",X"00",X"00",X"00",X"A0",X"46",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"D0",X"AA",X"9F",X"90",X"AD",X"AA",X"FF",X"9A",X"0A",X"AD",X"FF",X"FA",X"0A",X"A2",X"F3",X"FF",
		X"0A",X"FF",X"FB",X"FA",X"00",X"FF",X"FF",X"9A",X"00",X"FF",X"FF",X"AA",X"00",X"FB",X"FF",X"AA",
		X"FF",X"EF",X"FD",X"D0",X"FF",X"FF",X"A7",X"DD",X"FF",X"FB",X"7A",X"4D",X"3F",X"FF",X"90",X"42",
		X"FF",X"FF",X"80",X"A4",X"FF",X"00",X"00",X"A0",X"46",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"02",X"22",X"00",X"01",X"44",X"0B",X"2B",X"02",X"24",X"22",X"22",X"0E",X"40",X"32",X"B2",X"B3",
		X"0A",X"20",X"0B",X"B3",X"F2",X"D2",X"20",X"3E",X"FF",X"AA",X"D3",X"EE",X"BB",X"AA",X"A0",X"EE",
		X"DD",X"AA",X"AB",X"EF",X"DD",X"33",X"F2",X"DD",X"DD",X"AA",X"E2",X"DD",X"CE",X"DD",X"BB",X"DD",
		X"D0",X"DD",X"DD",X"DD",X"BB",X"00",X"DD",X"20",X"0A",X"BB",X"01",X"00",X"0A",X"0A",X"D2",X"D0",
		X"02",X"22",X"00",X"01",X"44",X"0B",X"2B",X"02",X"24",X"CC",X"22",X"0E",X"40",X"99",X"B2",X"B3",
		X"0A",X"11",X"0B",X"B3",X"F2",X"00",X"10",X"3E",X"FF",X"A0",X"CC",X"EE",X"BB",X"AA",X"A0",X"EE",
		X"DD",X"AA",X"AB",X"EF",X"DD",X"33",X"F2",X"DD",X"DD",X"AA",X"E2",X"DD",X"CE",X"DD",X"BB",X"DD",
		X"D0",X"DD",X"DD",X"DD",X"BB",X"00",X"DD",X"20",X"0A",X"BB",X"01",X"00",X"0A",X"0A",X"D2",X"D0",
		X"00",X"22",X"00",X"41",X"0B",X"0B",X"02",X"40",X"B2",X"BC",X"E0",X"00",X"22",X"11",X"BE",X"20",
		X"2D",X"91",X"AA",X"00",X"3B",X"99",X"AB",X"00",X"0D",X"99",X"32",X"00",X"90",X"AA",X"FF",X"D0",
		X"2B",X"AA",X"BB",X"DD",X"32",X"33",X"DD",X"ED",X"BD",X"E3",X"DD",X"0E",X"DD",X"DD",X"DD",X"BE",
		X"DF",X"DD",X"D0",X"EA",X"DD",X"0C",X"BB",X"A0",X"0C",X"BB",X"AA",X"70",X"22",X"BA",X"00",X"A6",
		X"00",X"07",X"77",X"77",X"00",X"07",X"FF",X"88",X"00",X"07",X"FF",X"88",X"00",X"07",X"FF",X"88",
		X"00",X"07",X"FF",X"88",X"00",X"07",X"FF",X"88",X"00",X"07",X"FF",X"88",X"00",X"07",X"FF",X"88",
		X"00",X"07",X"77",X"77",X"00",X"07",X"77",X"77",X"00",X"07",X"DD",X"DF",X"00",X"07",X"FD",X"FF",
		X"00",X"07",X"FD",X"DF",X"00",X"07",X"FD",X"FF",X"00",X"07",X"DD",X"FF",X"00",X"07",X"77",X"77",
		X"77",X"77",X"77",X"77",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"FF",X"FF",X"FF",X"DD",X"FF",X"FF",X"FF",X"DF",
		X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"DD",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"70",X"88",X"88",X"FF",X"70",X"88",X"88",X"FF",X"70",X"88",X"88",X"FF",X"70",
		X"88",X"88",X"FF",X"70",X"88",X"88",X"FF",X"70",X"88",X"88",X"FF",X"70",X"88",X"88",X"FF",X"70",
		X"77",X"77",X"77",X"70",X"77",X"77",X"77",X"70",X"DF",X"FF",X"FF",X"70",X"DF",X"FF",X"FF",X"70",
		X"DF",X"FF",X"FF",X"70",X"DF",X"FF",X"FF",X"70",X"DF",X"FF",X"FF",X"70",X"77",X"77",X"77",X"70",
		X"77",X"77",X"77",X"77",X"FF",X"88",X"88",X"88",X"FF",X"88",X"88",X"88",X"FF",X"88",X"88",X"88",
		X"FF",X"88",X"88",X"88",X"FF",X"88",X"88",X"88",X"FF",X"88",X"88",X"88",X"FF",X"88",X"88",X"88",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"FF",X"DD",X"DF",X"FF",X"FF",X"DF",X"FF",X"FF",
		X"FF",X"DD",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"DF",X"DF",X"DF",X"FF",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"FF",X"DF",X"DF",X"FF",X"FF",X"FF",X"DF",X"FF",
		X"FF",X"DF",X"DF",X"FF",X"FF",X"DF",X"DF",X"FF",X"FF",X"DF",X"DD",X"DF",X"77",X"77",X"77",X"77",
		X"77",X"77",X"00",X"00",X"8F",X"FF",X"00",X"00",X"8F",X"FF",X"00",X"00",X"8F",X"FF",X"00",X"00",
		X"8F",X"FF",X"00",X"00",X"8F",X"FF",X"00",X"00",X"8F",X"FF",X"00",X"00",X"8F",X"FF",X"00",X"00",
		X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"77",X"77",X"00",X"00",
		X"46",X"00",X"07",X"44",X"77",X"00",X"00",X"44",X"09",X"00",X"00",X"44",X"00",X"00",X"00",X"75",
		X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"31",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"13",X"00",X"00",X"11",X"11",X"00",
		X"46",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"02",X"11",
		X"00",X"00",X"07",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"72",
		X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"45",X"00",X"00",X"00",
		X"46",X"00",X"07",X"44",X"77",X"00",X"00",X"44",X"09",X"00",X"00",X"44",X"00",X"00",X"00",X"75",
		X"00",X"64",X"00",X"97",X"00",X"44",X"00",X"00",X"00",X"44",X"46",X"00",X"00",X"44",X"44",X"00",
		X"64",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"44",
		X"44",X"46",X"44",X"44",X"44",X"79",X"44",X"44",X"44",X"09",X"64",X"44",X"44",X"08",X"07",X"44",
		X"44",X"00",X"07",X"44",X"44",X"00",X"00",X"44",X"44",X"46",X"00",X"44",X"44",X"44",X"00",X"75",
		X"44",X"44",X"00",X"97",X"44",X"44",X"00",X"00",X"64",X"44",X"46",X"00",X"07",X"44",X"44",X"00",
		X"64",X"44",X"46",X"00",X"44",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"09",X"00",
		X"44",X"46",X"08",X"64",X"44",X"79",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"08",X"00",X"44",
		X"44",X"00",X"64",X"44",X"44",X"00",X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"77",X"64",X"44",X"44",X"00",X"07",X"44",X"44",X"00",
		X"07",X"44",X"46",X"00",X"09",X"44",X"77",X"00",X"00",X"64",X"09",X"00",X"00",X"07",X"00",X"00",
		X"00",X"07",X"00",X"64",X"00",X"09",X"00",X"44",X"60",X"00",X"00",X"44",X"45",X"00",X"00",X"44",
		X"46",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"64",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"46",X"00",X"00",X"44",X"44",X"00",
		X"64",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"44",
		X"44",X"46",X"44",X"44",X"44",X"79",X"44",X"44",X"44",X"09",X"64",X"44",X"44",X"08",X"07",X"44",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"46",X"00",X"00",X"44",X"44",X"00",X"00",
		X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"64",X"44",X"46",X"00",X"07",X"44",X"44",X"00",
		X"64",X"44",X"46",X"00",X"44",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"09",X"00",
		X"44",X"46",X"08",X"64",X"44",X"79",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"08",X"00",X"44",
		X"44",X"00",X"07",X"44",X"44",X"00",X"00",X"44",X"44",X"46",X"00",X"44",X"44",X"44",X"00",X"75",
		X"44",X"44",X"00",X"97",X"44",X"44",X"00",X"00",X"64",X"44",X"46",X"00",X"07",X"44",X"44",X"00",
		X"64",X"44",X"46",X"00",X"44",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"09",X"00",
		X"44",X"46",X"08",X"00",X"44",X"79",X"00",X"00",X"44",X"09",X"00",X"00",X"44",X"08",X"00",X"00",
		X"44",X"00",X"64",X"44",X"44",X"00",X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"77",X"64",X"44",X"44",X"00",X"07",X"44",X"44",X"00",
		X"07",X"44",X"46",X"00",X"09",X"44",X"77",X"00",X"00",X"64",X"09",X"00",X"00",X"07",X"00",X"00",
		X"00",X"07",X"00",X"64",X"00",X"09",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"46",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"44",X"60",X"00",X"00",X"44",X"45",X"00",X"00",X"44",
		X"46",X"00",X"07",X"44",X"77",X"00",X"00",X"44",X"09",X"00",X"00",X"44",X"00",X"00",X"00",X"75",
		X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"45",X"00",X"00",X"00",
		X"46",X"00",X"07",X"44",X"77",X"00",X"00",X"44",X"09",X"00",X"00",X"44",X"00",X"00",X"00",X"75",
		X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"44",X"60",X"00",X"00",X"44",X"45",X"00",X"00",X"44",
		X"46",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"45",X"00",X"00",X"00",
		X"00",X"00",X"07",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"75",
		X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"45",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"44",X"60",X"00",X"00",X"44",X"45",X"00",X"00",X"44",
		X"46",X"00",X"07",X"44",X"77",X"00",X"00",X"44",X"09",X"00",X"00",X"44",X"00",X"00",X"00",X"75",
		X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"46",X"00",X"64",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"64",X"44",X"46",X"00",X"44",X"44",X"77",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"64",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"44",
		X"44",X"46",X"44",X"44",X"44",X"79",X"44",X"44",X"44",X"09",X"64",X"44",X"44",X"08",X"07",X"44",
		X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"60",X"44",X"44",X"44",X"45",X"44",X"45",
		X"44",X"44",X"44",X"67",X"44",X"44",X"44",X"70",X"44",X"44",X"44",X"90",X"75",X"44",X"45",X"90",
		X"97",X"44",X"44",X"80",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"60",X"00",X"75",X"44",X"45",
		X"00",X"97",X"44",X"44",X"00",X"00",X"44",X"44",X"60",X"00",X"44",X"44",X"45",X"00",X"75",X"44",
		X"00",X"00",X"64",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"64",X"44",X"46",X"00",X"44",X"44",X"77",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"64",X"44",X"46",X"00",X"44",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"00",X"00",
		X"44",X"46",X"00",X"64",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"00",X"00",X"44",
		X"46",X"00",X"64",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"64",X"44",X"46",X"00",X"44",X"44",X"77",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"64",X"44",X"46",X"00",X"44",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"00",X"00",
		X"44",X"46",X"00",X"00",X"44",X"77",X"00",X"00",X"44",X"09",X"00",X"00",X"44",X"00",X"00",X"00",
		X"46",X"00",X"64",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"64",X"44",X"46",X"00",X"44",X"44",X"77",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"64",X"44",X"46",X"00",X"44",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"00",X"00",
		X"44",X"46",X"00",X"64",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"00",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"64",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"46",X"00",X"00",X"44",X"44",X"00",
		X"64",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"44",
		X"44",X"46",X"44",X"44",X"44",X"79",X"44",X"44",X"44",X"09",X"64",X"44",X"44",X"08",X"07",X"44",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"46",X"00",X"00",X"44",X"44",X"00",X"00",
		X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"64",X"44",X"46",X"00",X"07",X"44",X"44",X"00",
		X"64",X"44",X"46",X"00",X"44",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"09",X"00",
		X"44",X"46",X"08",X"00",X"44",X"79",X"00",X"00",X"44",X"09",X"00",X"00",X"44",X"08",X"00",X"00",
		X"44",X"00",X"64",X"44",X"44",X"00",X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"77",X"64",X"44",X"44",X"00",X"07",X"44",X"44",X"00",
		X"07",X"44",X"46",X"00",X"09",X"44",X"77",X"00",X"00",X"64",X"09",X"00",X"00",X"07",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"64",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"64",X"44",X"46",X"00",X"44",X"44",X"77",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"64",X"44",X"46",X"00",X"44",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"00",X"00",
		X"44",X"46",X"00",X"00",X"44",X"77",X"00",X"00",X"44",X"09",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"64",X"44",X"44",X"00",X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"77",X"64",X"44",X"44",X"90",X"07",X"44",X"44",X"90",
		X"64",X"44",X"44",X"80",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"44",
		X"44",X"46",X"44",X"44",X"44",X"97",X"44",X"44",X"44",X"90",X"64",X"44",X"44",X"80",X"07",X"44",
		X"00",X"00",X"64",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"64",X"44",X"46",X"00",X"44",X"44",X"77",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"64",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"44",
		X"44",X"46",X"44",X"44",X"44",X"79",X"44",X"44",X"44",X"09",X"64",X"44",X"44",X"08",X"07",X"44",
		X"44",X"00",X"64",X"44",X"44",X"00",X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"77",X"64",X"44",X"44",X"00",X"07",X"44",X"44",X"00",
		X"64",X"44",X"46",X"00",X"44",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"00",X"00",
		X"44",X"46",X"00",X"00",X"44",X"77",X"00",X"00",X"44",X"09",X"00",X"00",X"44",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"46",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"60",X"00",X"05",X"44",X"45",
		X"00",X"77",X"44",X"44",X"00",X"90",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"75",X"44",
		X"00",X"00",X"DC",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"DA",X"00",
		X"00",X"00",X"DA",X"00",X"00",X"00",X"DA",X"00",X"00",X"00",X"CA",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"DA",X"00",X"00",X"00",X"DA",X"00",X"00",X"00",X"DB",X"60",X"00",X"05",X"CB",X"45",
		X"00",X"77",X"CD",X"44",X"00",X"90",X"00",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"75",X"44",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"0F",X"00",X"00",X"0E",X"0F",X"00",X"00",X"0B",X"0F",X"00",
		X"00",X"0B",X"0F",X"00",X"00",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"00",X"00",X"0F",X"FC",X"00",
		X"00",X"0F",X"CC",X"00",X"00",X"0F",X"CE",X"00",X"00",X"0B",X"CF",X"00",X"00",X"00",X"DF",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"EC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"30",X"00",X"00",X"11",X"12",X"00",X"00",
		X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"30",X"00",X"72",X"11",X"12",X"00",
		X"DD",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CD",X"00",X"00",X"00",X"CD",X"00",X"00",X"00",
		X"CD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",
		X"CD",X"00",X"00",X"00",X"CD",X"00",X"00",X"00",X"CD",X"30",X"00",X"00",X"DC",X"02",X"00",X"00",
		X"BC",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"11",X"11",X"30",X"00",X"72",X"11",X"12",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"CD",X"00",X"00",X"00",
		X"ED",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"2D",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"C2",X"00",X"00",X"0D",X"D3",
		X"00",X"00",X"0D",X"DB",X"00",X"00",X"0B",X"DD",X"00",X"00",X"03",X"3D",X"00",X"00",X"03",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",
		X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"3D",X"00",X"00",X"00",X"2C",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"0D",X"00",X"D0",X"0D",X"0D",X"00",X"D0",X"0C",X"00",X"00",X"00",X"0C",X"00",
		X"00",X"00",X"0D",X"DF",X"00",X"00",X"0D",X"DF",X"00",X"00",X"00",X"3D",X"00",X"00",X"00",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"CD",
		X"00",X"00",X"00",X"3D",X"00",X"00",X"00",X"0D",X"00",X"00",X"0D",X"0D",X"00",X"00",X"03",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"D0",
		X"00",X"00",X"0C",X"3F",X"00",X"00",X"0C",X"2D",X"00",X"00",X"0B",X"D2",X"D0",X"00",X"0C",X"D3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"CD",
		X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"D0",X"00",X"00",X"0D",X"30",X"00",X"00",X"0D",X"2D",X"00",X"00",X"0C",X"D2",
		X"00",X"D0",X"0C",X"D3",X"B0",X"D0",X"0C",X"DD",X"D0",X"D0",X"0C",X"DD",X"00",X"00",X"0B",X"DF",
		X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",
		X"00",X"00",X"0D",X"30",X"00",X"00",X"D0",X"2D",X"00",X"D0",X"D0",X"D2",X"00",X"D0",X"DD",X"D3",
		X"0D",X"D0",X"03",X"DD",X"00",X"D0",X"03",X"DD",X"00",X"D0",X"03",X"DD",X"00",X"00",X"02",X"3F",
		X"00",X"00",X"6C",X"CF",X"D0",X"00",X"FC",X"FF",X"B0",X"00",X"FD",X"FF",X"C0",X"00",X"FD",X"FF",
		X"00",X"DF",X"DF",X"F6",X"00",X"BF",X"FF",X"77",X"00",X"CF",X"FF",X"00",X"D0",X"DD",X"FF",X"00",
		X"DF",X"CF",X"F4",X"00",X"DD",X"FF",X"44",X"00",X"CD",X"FF",X"44",X"46",X"3D",X"FF",X"44",X"44",
		X"3F",X"F6",X"44",X"44",X"FF",X"79",X"44",X"44",X"FF",X"09",X"64",X"44",X"FF",X"08",X"07",X"44",
		X"00",X"00",X"6D",X"CF",X"30",X"00",X"FD",X"FF",X"30",X"00",X"FB",X"FF",X"C0",X"00",X"DF",X"FF",
		X"D0",X"DF",X"DF",X"F6",X"00",X"DF",X"FF",X"77",X"00",X"DD",X"FF",X"00",X"D0",X"DD",X"FF",X"00",
		X"BD",X"CF",X"F4",X"00",X"3D",X"FF",X"44",X"00",X"33",X"FF",X"44",X"46",X"D2",X"FF",X"44",X"44",
		X"DF",X"F6",X"44",X"44",X"FF",X"79",X"44",X"44",X"FF",X"09",X"64",X"44",X"FF",X"08",X"07",X"44",
		X"D0",X"00",X"6D",X"CF",X"D0",X"00",X"FC",X"FF",X"00",X"00",X"D3",X"FF",X"00",X"00",X"DF",X"FF",
		X"00",X"6F",X"DF",X"F6",X"00",X"DF",X"FF",X"77",X"00",X"DD",X"FF",X"00",X"D0",X"CD",X"FF",X"00",
		X"3D",X"CF",X"F4",X"00",X"2C",X"FF",X"44",X"00",X"23",X"FF",X"44",X"46",X"D2",X"FF",X"44",X"44",
		X"DF",X"F6",X"44",X"44",X"FF",X"79",X"44",X"44",X"FF",X"09",X"64",X"44",X"FF",X"08",X"07",X"44",
		X"00",X"00",X"62",X"DF",X"0D",X"00",X"F2",X"FF",X"D0",X"00",X"D3",X"FF",X"D0",X"00",X"DD",X"FF",
		X"00",X"DF",X"DF",X"F6",X"00",X"3F",X"FF",X"77",X"30",X"2D",X"FF",X"00",X"2B",X"CD",X"FF",X"00",
		X"B3",X"DF",X"F4",X"00",X"D2",X"FF",X"44",X"00",X"DC",X"FF",X"44",X"46",X"DD",X"FF",X"44",X"44",
		X"DF",X"F6",X"44",X"44",X"FF",X"79",X"44",X"44",X"FF",X"09",X"64",X"44",X"FF",X"08",X"07",X"44",
		X"00",X"00",X"63",X"3F",X"D0",X"00",X"FD",X"FF",X"D0",X"00",X"DD",X"FF",X"C0",X"00",X"DD",X"FF",
		X"30",X"BF",X"DF",X"F6",X"2C",X"2F",X"FF",X"77",X"3C",X"3C",X"FF",X"00",X"B3",X"BD",X"FF",X"00",
		X"C3",X"DF",X"F4",X"00",X"DB",X"FF",X"44",X"00",X"DC",X"FF",X"44",X"46",X"DD",X"FF",X"44",X"44",
		X"2F",X"F6",X"44",X"44",X"FF",X"79",X"44",X"44",X"FF",X"09",X"64",X"44",X"FF",X"08",X"07",X"44",
		X"00",X"00",X"6C",X"CF",X"D0",X"00",X"FC",X"FF",X"B0",X"00",X"FD",X"FF",X"C0",X"00",X"FD",X"FF",
		X"00",X"DF",X"DF",X"F6",X"00",X"BF",X"FF",X"77",X"00",X"CF",X"FF",X"00",X"D0",X"DD",X"FF",X"00",
		X"DF",X"CF",X"FF",X"00",X"DD",X"FF",X"FF",X"00",X"CD",X"FF",X"FF",X"F6",X"3D",X"FF",X"FF",X"FF",
		X"3F",X"F6",X"FF",X"FF",X"FF",X"79",X"FF",X"FF",X"FF",X"09",X"6F",X"FF",X"FF",X"08",X"07",X"FF",
		X"00",X"00",X"6D",X"CF",X"30",X"00",X"FD",X"FF",X"30",X"00",X"FB",X"FF",X"C0",X"00",X"DF",X"FF",
		X"D0",X"DF",X"DF",X"F6",X"00",X"DF",X"FF",X"77",X"00",X"DD",X"FF",X"00",X"D0",X"DD",X"FF",X"00",
		X"BD",X"CF",X"FF",X"00",X"3D",X"FF",X"FF",X"00",X"33",X"FF",X"FF",X"F6",X"D2",X"FF",X"FF",X"FF",
		X"DF",X"F6",X"FF",X"FF",X"FF",X"79",X"FF",X"FF",X"FF",X"09",X"6F",X"FF",X"FF",X"08",X"07",X"FF",
		X"D0",X"00",X"6D",X"CF",X"D0",X"00",X"FC",X"FF",X"00",X"00",X"D3",X"FF",X"00",X"00",X"DF",X"FF",
		X"00",X"6F",X"DF",X"F6",X"00",X"DF",X"FF",X"77",X"00",X"DD",X"FF",X"00",X"D0",X"CD",X"FF",X"00",
		X"3D",X"CF",X"FF",X"00",X"2C",X"FF",X"FF",X"00",X"23",X"FF",X"FF",X"F6",X"D2",X"FF",X"FF",X"FF",
		X"DF",X"F6",X"FF",X"FF",X"FF",X"79",X"FF",X"FF",X"FF",X"09",X"6F",X"FF",X"FF",X"08",X"07",X"FF",
		X"00",X"00",X"62",X"DF",X"0D",X"00",X"F2",X"FF",X"D0",X"00",X"D3",X"FF",X"D0",X"00",X"DD",X"FF",
		X"00",X"DF",X"DF",X"F6",X"00",X"3F",X"FF",X"77",X"30",X"2D",X"FF",X"00",X"2B",X"CD",X"FF",X"00",
		X"B3",X"DF",X"FF",X"00",X"D2",X"FF",X"FF",X"00",X"DC",X"FF",X"FF",X"F6",X"DD",X"FF",X"FF",X"FF",
		X"DF",X"F6",X"FF",X"FF",X"FF",X"79",X"FF",X"FF",X"FF",X"09",X"6F",X"FF",X"FF",X"08",X"07",X"FF",
		X"00",X"00",X"63",X"3F",X"D0",X"00",X"FD",X"FF",X"D0",X"00",X"DD",X"FF",X"C0",X"00",X"DD",X"FF",
		X"30",X"BF",X"DF",X"F6",X"2C",X"2F",X"FF",X"77",X"3C",X"3C",X"FF",X"00",X"B3",X"BD",X"FF",X"00",
		X"C3",X"DF",X"FF",X"00",X"DB",X"FF",X"FF",X"00",X"DC",X"FF",X"FF",X"F6",X"DD",X"FF",X"FF",X"FF",
		X"2F",X"F6",X"FF",X"FF",X"FF",X"79",X"FF",X"FF",X"FF",X"09",X"6F",X"FF",X"FF",X"08",X"07",X"FF",
		X"00",X"00",X"6C",X"CF",X"D0",X"00",X"FC",X"FF",X"B0",X"00",X"FD",X"FF",X"C0",X"00",X"FD",X"FF",
		X"00",X"DF",X"DF",X"F6",X"00",X"BF",X"FF",X"77",X"00",X"CF",X"FF",X"D0",X"D0",X"DD",X"FF",X"C0",
		X"DF",X"CF",X"FF",X"2D",X"DD",X"FF",X"FF",X"23",X"CD",X"FF",X"FF",X"C2",X"3D",X"FF",X"FD",X"D3",
		X"3F",X"F6",X"FD",X"DB",X"FF",X"79",X"FB",X"DD",X"FF",X"09",X"63",X"3D",X"FF",X"08",X"03",X"2D",
		X"00",X"00",X"6D",X"CF",X"30",X"00",X"FD",X"FF",X"30",X"00",X"FB",X"FF",X"C0",X"00",X"DF",X"DF",
		X"D0",X"DF",X"DF",X"D6",X"00",X"DF",X"FF",X"3D",X"00",X"DD",X"FF",X"2C",X"D0",X"DD",X"FF",X"03",
		X"BD",X"CF",X"FF",X"0D",X"3D",X"DF",X"FD",X"0D",X"33",X"DF",X"FC",X"F6",X"D2",X"FF",X"FC",X"FF",
		X"DF",X"F6",X"FD",X"DF",X"FF",X"79",X"FD",X"DF",X"FF",X"09",X"6F",X"3D",X"FF",X"08",X"07",X"2D",
		X"D0",X"00",X"6D",X"CF",X"D0",X"00",X"FC",X"DF",X"00",X"00",X"D3",X"DF",X"00",X"00",X"DF",X"CD",
		X"00",X"6F",X"DF",X"3D",X"00",X"DF",X"FF",X"7D",X"00",X"DD",X"FD",X"0D",X"D0",X"CD",X"F3",X"00",
		X"3D",X"CF",X"FB",X"00",X"2C",X"FF",X"FF",X"00",X"23",X"FF",X"FF",X"F6",X"D2",X"FF",X"FC",X"DF",
		X"DF",X"F6",X"FC",X"3F",X"FF",X"79",X"FC",X"2D",X"FF",X"09",X"6B",X"D2",X"DF",X"08",X"0C",X"D3",
		X"00",X"00",X"62",X"DF",X"0D",X"00",X"F2",X"DF",X"D0",X"00",X"D3",X"DF",X"D0",X"00",X"DD",X"CD",
		X"00",X"DF",X"DF",X"FD",X"00",X"3F",X"FF",X"77",X"30",X"2D",X"FF",X"00",X"2B",X"CD",X"FF",X"00",
		X"B3",X"DF",X"FF",X"D0",X"D2",X"FF",X"FD",X"30",X"DC",X"FF",X"FD",X"2D",X"DD",X"FF",X"FC",X"D2",
		X"DF",X"D6",X"FC",X"D3",X"BF",X"D9",X"FC",X"DD",X"DF",X"D9",X"6C",X"DD",X"FF",X"08",X"0B",X"DF",
		X"00",X"00",X"63",X"DF",X"D0",X"00",X"FD",X"DF",X"D0",X"00",X"DD",X"FF",X"C0",X"00",X"DD",X"FF",
		X"30",X"BF",X"DF",X"F6",X"2C",X"2F",X"FF",X"77",X"3C",X"3C",X"FF",X"00",X"B3",X"BD",X"FF",X"D0",
		X"C3",X"DF",X"FD",X"30",X"DB",X"FF",X"DF",X"2D",X"DC",X"DF",X"DF",X"D2",X"DD",X"DF",X"DD",X"D3",
		X"2D",X"D6",X"F3",X"DD",X"FF",X"D9",X"F3",X"DD",X"FF",X"D9",X"63",X"DD",X"FF",X"08",X"02",X"3F",
		X"FF",X"00",X"6C",X"CF",X"DF",X"00",X"FC",X"FF",X"BF",X"F6",X"FD",X"FF",X"CF",X"FF",X"FD",X"FF",
		X"FF",X"DF",X"DF",X"F6",X"FF",X"BF",X"FF",X"77",X"6F",X"CF",X"FF",X"90",X"D7",X"DD",X"FF",X"90",
		X"DF",X"CF",X"F4",X"80",X"DD",X"FF",X"44",X"00",X"CD",X"FF",X"44",X"46",X"3D",X"FF",X"44",X"44",
		X"3F",X"F6",X"44",X"44",X"FF",X"97",X"44",X"44",X"FF",X"90",X"64",X"44",X"FF",X"80",X"07",X"44",
		X"FF",X"00",X"6D",X"CF",X"3F",X"00",X"FD",X"FF",X"3F",X"F6",X"FB",X"FF",X"CF",X"FF",X"DF",X"FF",
		X"DF",X"DF",X"DF",X"F6",X"FF",X"DF",X"FF",X"77",X"6F",X"DD",X"FF",X"90",X"D7",X"DD",X"FF",X"90",
		X"BD",X"CF",X"F4",X"80",X"3D",X"FF",X"44",X"00",X"33",X"FF",X"44",X"46",X"D2",X"FF",X"44",X"44",
		X"DF",X"F6",X"44",X"44",X"FF",X"97",X"44",X"44",X"FF",X"90",X"64",X"44",X"FF",X"80",X"07",X"44",
		X"DF",X"00",X"6D",X"CF",X"DF",X"00",X"FC",X"FF",X"FF",X"F6",X"D3",X"FF",X"FF",X"FF",X"DF",X"FF",
		X"FF",X"FF",X"DF",X"F6",X"FF",X"DF",X"FF",X"77",X"6F",X"DD",X"FF",X"90",X"D7",X"CD",X"FF",X"90",
		X"3D",X"CF",X"F4",X"80",X"2C",X"FF",X"44",X"00",X"23",X"FF",X"44",X"46",X"D2",X"FF",X"44",X"44",
		X"DF",X"F6",X"44",X"44",X"FF",X"97",X"44",X"44",X"FF",X"90",X"64",X"44",X"FF",X"80",X"07",X"44",
		X"FF",X"00",X"62",X"DF",X"FD",X"00",X"F2",X"FF",X"DF",X"F6",X"D3",X"FF",X"DF",X"FF",X"DD",X"FF",
		X"FF",X"DF",X"DF",X"F6",X"FF",X"3F",X"FF",X"77",X"3F",X"2D",X"FF",X"90",X"2B",X"CD",X"FF",X"90",
		X"B3",X"DF",X"F4",X"80",X"D2",X"FF",X"44",X"00",X"DC",X"FF",X"44",X"46",X"DD",X"FF",X"44",X"44",
		X"DF",X"F6",X"44",X"44",X"FF",X"97",X"44",X"44",X"FF",X"90",X"64",X"44",X"FF",X"80",X"07",X"44",
		X"FF",X"00",X"63",X"3F",X"DF",X"00",X"FD",X"FF",X"DF",X"F6",X"DD",X"FF",X"CF",X"FF",X"DD",X"FF",
		X"3F",X"BF",X"DF",X"F6",X"2C",X"2F",X"FF",X"77",X"3C",X"3C",X"FF",X"90",X"B3",X"BD",X"FF",X"90",
		X"C3",X"DF",X"F4",X"80",X"DB",X"FF",X"44",X"00",X"DC",X"FF",X"44",X"46",X"DD",X"FF",X"44",X"44",
		X"2F",X"F6",X"44",X"44",X"FF",X"97",X"44",X"44",X"FF",X"90",X"64",X"44",X"FF",X"80",X"07",X"44",
		X"FF",X"00",X"6C",X"CF",X"DF",X"00",X"FC",X"FF",X"BF",X"F6",X"FD",X"FF",X"CF",X"FF",X"FD",X"FF",
		X"FF",X"DF",X"DF",X"F6",X"FF",X"BF",X"FF",X"77",X"6F",X"CF",X"FF",X"90",X"D7",X"DD",X"FF",X"90",
		X"DF",X"CF",X"FF",X"80",X"DD",X"FF",X"FF",X"00",X"CD",X"FF",X"FF",X"F6",X"3D",X"FF",X"FF",X"FF",
		X"3F",X"F6",X"FF",X"FF",X"FF",X"97",X"FF",X"FF",X"FF",X"90",X"6F",X"FF",X"FF",X"80",X"07",X"FF",
		X"FF",X"00",X"6D",X"CF",X"3F",X"00",X"FD",X"FF",X"3F",X"F6",X"FB",X"FF",X"CF",X"FF",X"DF",X"FF",
		X"DF",X"DF",X"DF",X"F6",X"FF",X"DF",X"FF",X"77",X"6F",X"DD",X"FF",X"90",X"D7",X"DD",X"FF",X"90",
		X"BD",X"CF",X"FF",X"80",X"3D",X"FF",X"FF",X"00",X"33",X"FF",X"FF",X"F6",X"D2",X"FF",X"FF",X"FF",
		X"DF",X"F6",X"FF",X"FF",X"FF",X"97",X"FF",X"FF",X"FF",X"90",X"6F",X"FF",X"FF",X"80",X"07",X"FF",
		X"DF",X"00",X"6D",X"CF",X"DF",X"00",X"FC",X"FF",X"FF",X"F6",X"D3",X"FF",X"FF",X"FF",X"DF",X"FF",
		X"FF",X"FF",X"DF",X"F6",X"FF",X"DF",X"FF",X"77",X"6F",X"DD",X"FF",X"90",X"D7",X"CD",X"FF",X"90",
		X"3D",X"CF",X"FF",X"80",X"2C",X"FF",X"FF",X"00",X"23",X"FF",X"FF",X"F6",X"D2",X"FF",X"FF",X"FF",
		X"DF",X"F6",X"FF",X"FF",X"FF",X"97",X"FF",X"FF",X"FF",X"90",X"6F",X"FF",X"FF",X"80",X"07",X"FF",
		X"FF",X"00",X"62",X"DF",X"FD",X"00",X"F2",X"FF",X"DF",X"F6",X"D3",X"FF",X"DF",X"FF",X"DD",X"FF",
		X"FF",X"DF",X"DF",X"F6",X"FF",X"3F",X"FF",X"77",X"3F",X"2D",X"FF",X"90",X"2B",X"CD",X"FF",X"90",
		X"B3",X"DF",X"FF",X"80",X"D2",X"FF",X"FF",X"00",X"DC",X"FF",X"FF",X"F6",X"DD",X"FF",X"FF",X"FF",
		X"DF",X"F6",X"FF",X"FF",X"FF",X"97",X"FF",X"FF",X"FF",X"90",X"6F",X"FF",X"FF",X"80",X"07",X"FF",
		X"FF",X"00",X"63",X"3F",X"DF",X"00",X"FD",X"FF",X"DF",X"F6",X"DD",X"FF",X"CF",X"FF",X"DD",X"FF",
		X"3F",X"BF",X"DF",X"F6",X"2C",X"2F",X"FF",X"77",X"3C",X"3C",X"FF",X"90",X"B3",X"BD",X"FF",X"90",
		X"C3",X"DF",X"FF",X"80",X"DB",X"FF",X"FF",X"00",X"DC",X"FF",X"FF",X"F6",X"DD",X"FF",X"FF",X"FF",
		X"2F",X"F6",X"FF",X"FF",X"FF",X"97",X"FF",X"FF",X"FF",X"90",X"6F",X"FF",X"FF",X"80",X"07",X"FF",
		X"FF",X"00",X"6C",X"CF",X"DF",X"00",X"FC",X"FF",X"BF",X"F6",X"FD",X"FF",X"CF",X"FF",X"FD",X"FF",
		X"FF",X"DF",X"DF",X"F6",X"FF",X"BF",X"FF",X"77",X"6F",X"CF",X"FF",X"D0",X"D7",X"DD",X"FF",X"C0",
		X"DF",X"CF",X"FF",X"2D",X"DD",X"FF",X"FF",X"23",X"CD",X"FF",X"FF",X"C2",X"3D",X"FF",X"FD",X"D3",
		X"3F",X"F6",X"FD",X"DB",X"FF",X"97",X"FB",X"DD",X"FF",X"90",X"63",X"3D",X"FF",X"80",X"03",X"2D",
		X"FF",X"00",X"6D",X"CF",X"3F",X"00",X"FD",X"FF",X"3F",X"F6",X"FB",X"FF",X"CF",X"FF",X"DF",X"DF",
		X"DF",X"DF",X"DF",X"D6",X"FF",X"DF",X"FF",X"3D",X"6F",X"DD",X"FF",X"2C",X"D7",X"DD",X"FF",X"93",
		X"BD",X"CF",X"FF",X"8D",X"3D",X"DF",X"FD",X"0D",X"33",X"DF",X"FC",X"F6",X"D2",X"FF",X"FC",X"FF",
		X"DF",X"F6",X"FD",X"DF",X"FF",X"97",X"FD",X"DF",X"FF",X"90",X"6F",X"3D",X"FF",X"80",X"07",X"2D",
		X"DF",X"00",X"6D",X"CF",X"DF",X"00",X"FC",X"DF",X"FF",X"F6",X"D3",X"DF",X"FF",X"FF",X"DF",X"CD",
		X"FF",X"FF",X"DF",X"3D",X"FF",X"DF",X"FF",X"7D",X"6F",X"DD",X"FD",X"9D",X"D7",X"CD",X"F3",X"90",
		X"3D",X"CF",X"FB",X"80",X"2C",X"FF",X"FF",X"00",X"23",X"FF",X"FF",X"F6",X"D2",X"FF",X"FC",X"DF",
		X"DF",X"F6",X"FC",X"3F",X"FF",X"97",X"FC",X"2D",X"FF",X"90",X"6B",X"D2",X"DF",X"80",X"0C",X"D3",
		X"FF",X"00",X"62",X"DF",X"FD",X"00",X"F2",X"DF",X"DF",X"F6",X"D3",X"DF",X"DF",X"FF",X"DD",X"CD",
		X"FF",X"DF",X"DF",X"FD",X"FF",X"3F",X"FF",X"77",X"3F",X"2D",X"FF",X"90",X"2B",X"CD",X"FF",X"90",
		X"B3",X"DF",X"FF",X"D0",X"D2",X"FF",X"FD",X"30",X"DC",X"FF",X"FD",X"2D",X"DD",X"FF",X"FC",X"D2",
		X"DF",X"D6",X"FC",X"D3",X"BF",X"D7",X"FC",X"DD",X"DF",X"D0",X"6C",X"DD",X"FF",X"80",X"0B",X"DF",
		X"FF",X"00",X"63",X"DF",X"DF",X"00",X"FD",X"DF",X"DF",X"F6",X"DD",X"FF",X"CF",X"FF",X"DD",X"FF",
		X"3F",X"BF",X"DF",X"F6",X"2C",X"2F",X"FF",X"77",X"3C",X"3C",X"FF",X"90",X"B3",X"BD",X"FF",X"D0",
		X"C3",X"DF",X"FD",X"30",X"DB",X"FF",X"DF",X"2D",X"DC",X"DF",X"DF",X"D2",X"DD",X"DF",X"DD",X"D3",
		X"2D",X"D6",X"F3",X"DD",X"FF",X"D7",X"F3",X"DD",X"FF",X"D0",X"63",X"DD",X"FF",X"80",X"02",X"3F",
		X"00",X"00",X"6F",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"6F",X"FF",X"F6",X"00",X"FF",X"FF",X"77",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"6F",X"FF",X"F4",X"00",X"FF",X"FF",X"44",X"00",X"FF",X"FF",X"44",X"46",X"FF",X"FF",X"44",X"44",
		X"FF",X"F6",X"44",X"44",X"FF",X"79",X"44",X"44",X"FF",X"09",X"64",X"44",X"FF",X"08",X"07",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"6F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"07",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"75",
		X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"6F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"07",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"75",
		X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"F4",X"00",X"64",X"44",X"44",X"00",X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"77",X"64",X"44",X"44",X"90",X"07",X"44",X"44",X"90",
		X"64",X"44",X"44",X"80",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"46",X"44",X"44",X"44",X"44",
		X"44",X"46",X"44",X"44",X"44",X"97",X"44",X"44",X"44",X"90",X"64",X"44",X"44",X"80",X"07",X"44",
		X"FF",X"00",X"6F",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"77",X"6F",X"FF",X"FF",X"90",X"07",X"FF",X"FF",X"90",
		X"6F",X"FF",X"F4",X"80",X"FF",X"FF",X"44",X"00",X"FF",X"FF",X"44",X"46",X"FF",X"FF",X"44",X"44",
		X"FF",X"F6",X"44",X"44",X"FF",X"97",X"44",X"44",X"FF",X"90",X"64",X"44",X"FF",X"80",X"07",X"44",
		X"FF",X"00",X"6F",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"77",X"6F",X"FF",X"FF",X"90",X"07",X"FF",X"FF",X"90",
		X"6F",X"FF",X"FF",X"80",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F6",X"FF",X"FF",X"FF",X"97",X"FF",X"FF",X"FF",X"90",X"6F",X"FF",X"FF",X"80",X"07",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
