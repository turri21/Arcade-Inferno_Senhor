library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity inferno_prog2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)

	-- signals that carry the ROM data from the MiSTer disk
	--dn_addr : in  std_logic_vector(15 downto 0);
	--dn_dout : in  std_logic_vector(7 downto 0);
	--dn_wr   : in  std_logic
);
end entity;

architecture prom of inferno_prog2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	
	signal rom_data: rom := (
		X"1A",X"F0",X"10",X"CE",X"BF",X"60",X"7E",X"E0",X"B6",X"BD",X"E9",X"E4",X"49",X"00",X"05",X"39",
		X"BD",X"E9",X"E4",X"49",X"03",X"05",X"39",X"BD",X"E9",X"E4",X"49",X"06",X"05",X"39",X"BD",X"E9",
		X"E4",X"49",X"09",X"05",X"39",X"BD",X"E9",X"E4",X"49",X"0C",X"05",X"39",X"BD",X"E9",X"E4",X"49",
		X"0F",X"05",X"39",X"BD",X"E9",X"E4",X"49",X"12",X"05",X"39",X"BD",X"E9",X"E4",X"49",X"15",X"05",
		X"39",X"BD",X"E9",X"E4",X"49",X"18",X"05",X"39",X"BD",X"E9",X"E4",X"49",X"1B",X"05",X"39",X"BD",
		X"E9",X"E4",X"49",X"1E",X"05",X"39",X"BD",X"E9",X"E4",X"49",X"21",X"05",X"39",X"7E",X"EA",X"90",
		X"7E",X"EA",X"B1",X"7E",X"E4",X"5C",X"7E",X"E4",X"37",X"7E",X"E3",X"B5",X"7E",X"E3",X"48",X"7E",
		X"E7",X"23",X"7E",X"E7",X"46",X"7E",X"E7",X"62",X"7E",X"E4",X"5E",X"EB",X"2A",X"7E",X"E3",X"46",
		X"7E",X"E4",X"8D",X"7E",X"E5",X"A5",X"E7",X"0B",X"7E",X"E4",X"C7",X"7E",X"E5",X"0B",X"E4",X"8C",
		X"7E",X"E5",X"6D",X"7E",X"E8",X"22",X"7E",X"E5",X"8B",X"7E",X"E9",X"E4",X"EA",X"13",X"7E",X"E7",
		X"93",X"7E",X"E7",X"7E",X"7E",X"E7",X"F3",X"7E",X"E7",X"A8",X"7E",X"E3",X"5B",X"7E",X"E4",X"BF",
		X"7E",X"E4",X"A5",X"7E",X"EA",X"F1",X"86",X"90",X"1F",X"8B",X"7F",X"BF",X"FF",X"7F",X"C8",X"00",
		X"86",X"C0",X"B7",X"C9",X"8C",X"8E",X"00",X"00",X"1F",X"13",X"86",X"14",X"B7",X"C9",X"00",X"EF",
		X"81",X"8C",X"BF",X"80",X"25",X"F6",X"8E",X"D0",X"00",X"B7",X"C9",X"00",X"EF",X"81",X"8C",X"DF",
		X"FF",X"25",X"F6",X"C6",X"03",X"F7",X"BF",X"FF",X"F7",X"C8",X"00",X"10",X"8E",X"00",X"00",X"8E",
		X"80",X"00",X"B7",X"C9",X"00",X"10",X"AF",X"89",X"40",X"00",X"EF",X"81",X"10",X"AF",X"89",X"40",
		X"00",X"EF",X"81",X"8C",X"87",X"FF",X"25",X"EA",X"CC",X"00",X"01",X"F7",X"BF",X"FF",X"F7",X"C8",
		X"00",X"B7",X"C9",X"81",X"B7",X"C9",X"83",X"B7",X"C9",X"85",X"B7",X"C9",X"87",X"C6",X"35",X"FD",
		X"C9",X"80",X"C6",X"34",X"FD",X"C9",X"84",X"FD",X"C9",X"86",X"43",X"C6",X"2C",X"FD",X"C9",X"82",
		X"BD",X"E7",X"7E",X"7F",X"CB",X"C0",X"CE",X"D1",X"2F",X"DF",X"00",X"86",X"10",X"30",X"C8",X"6F",
		X"AF",X"C4",X"33",X"88",X"6F",X"EF",X"84",X"4A",X"26",X"F3",X"4F",X"5F",X"ED",X"84",X"0A",X"05",
		X"86",X"07",X"B7",X"CB",X"00",X"4C",X"B7",X"CB",X"20",X"8E",X"EB",X"2A",X"BD",X"E7",X"23",X"86",
		X"01",X"B7",X"CB",X"A0",X"7F",X"CB",X"80",X"86",X"0A",X"B7",X"CB",X"40",X"7F",X"CB",X"60",X"CC",
		X"0E",X"10",X"DD",X"6B",X"8E",X"CD",X"00",X"BD",X"00",X"27",X"1F",X"98",X"81",X"20",X"22",X"06",
		X"84",X"0F",X"81",X"09",X"23",X"07",X"5F",X"8E",X"CD",X"00",X"BD",X"00",X"30",X"D7",X"E1",X"CE",
		X"90",X"02",X"10",X"8E",X"11",X"00",X"4F",X"5F",X"BD",X"E4",X"5E",X"8E",X"90",X"14",X"9F",X"0E",
		X"0C",X"13",X"1C",X"EF",X"DE",X"04",X"2A",X"04",X"AE",X"56",X"2B",X"03",X"7E",X"E1",X"D3",X"10",
		X"8E",X"90",X"0E",X"A6",X"48",X"A0",X"08",X"25",X"12",X"22",X"06",X"A6",X"42",X"A1",X"02",X"22",
		X"0A",X"EC",X"16",X"AF",X"36",X"EF",X"16",X"ED",X"56",X"1E",X"13",X"31",X"C4",X"33",X"84",X"AE",
		X"16",X"2B",X"E0",X"86",X"05",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"DE",X"04",X"DF",X"0A",X"DF",
		X"08",X"CC",X"B7",X"89",X"FD",X"B8",X"27",X"10",X"8E",X"B8",X"AB",X"10",X"9F",X"16",X"DE",X"0A",
		X"2A",X"0D",X"A6",X"5E",X"81",X"40",X"24",X"07",X"AD",X"D8",X"F8",X"EE",X"56",X"2B",X"F3",X"DF",
		X"0A",X"6F",X"A0",X"10",X"9F",X"18",X"DE",X"0A",X"2A",X"0D",X"A6",X"5E",X"2B",X"07",X"AD",X"D8",
		X"F8",X"EE",X"56",X"2B",X"F5",X"DF",X"0A",X"86",X"60",X"BD",X"E3",X"79",X"DE",X"08",X"2A",X"0F",
		X"A6",X"5E",X"81",X"40",X"24",X"07",X"AD",X"D8",X"5A",X"EE",X"56",X"2B",X"F3",X"DF",X"08",X"6F",
		X"A0",X"10",X"9F",X"1A",X"DE",X"0A",X"2A",X"0F",X"A6",X"5E",X"81",X"C0",X"24",X"07",X"AD",X"D8",
		X"F8",X"EE",X"56",X"2B",X"F3",X"DF",X"0A",X"86",X"A0",X"BD",X"E3",X"79",X"DE",X"08",X"2A",X"0D",
		X"A6",X"5E",X"2B",X"07",X"AD",X"D8",X"5A",X"EE",X"56",X"2B",X"F5",X"DF",X"08",X"6F",X"A0",X"10",
		X"9F",X"1C",X"DE",X"0A",X"2A",X"07",X"AD",X"D8",X"F8",X"EE",X"56",X"2B",X"F9",X"86",X"FF",X"BD",
		X"E3",X"79",X"DE",X"08",X"2A",X"07",X"AD",X"D8",X"5A",X"EE",X"56",X"2B",X"F9",X"6F",X"A0",X"0F",
		X"13",X"86",X"01",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"1A",X"10",X"D6",X"4F",X"0F",X"4F",X"1C",
		X"EF",X"C4",X"38",X"27",X"03",X"BD",X"11",X"3B",X"96",X"4B",X"27",X"28",X"0A",X"4B",X"26",X"63",
		X"9E",X"4D",X"27",X"20",X"EC",X"81",X"2B",X"03",X"8E",X"00",X"00",X"9F",X"4D",X"D7",X"4B",X"84",
		X"7F",X"97",X"B6",X"8E",X"E7",X"B6",X"1F",X"89",X"3A",X"81",X"01",X"27",X"46",X"A6",X"84",X"B7",
		X"C9",X"82",X"20",X"3F",X"DC",X"A7",X"91",X"A9",X"22",X"02",X"DC",X"A9",X"91",X"AB",X"22",X"02",
		X"DC",X"AB",X"91",X"AD",X"22",X"02",X"DC",X"AD",X"91",X"AF",X"22",X"02",X"DC",X"AF",X"91",X"B1",
		X"22",X"02",X"DC",X"B1",X"91",X"B3",X"22",X"02",X"DC",X"B3",X"97",X"4C",X"D1",X"B6",X"27",X"13",
		X"D7",X"B6",X"C1",X"35",X"26",X"04",X"86",X"36",X"97",X"B0",X"8E",X"E7",X"B6",X"3A",X"E6",X"84",
		X"F7",X"C9",X"82",X"CE",X"90",X"02",X"DF",X"21",X"CC",X"E3",X"11",X"DD",X"73",X"10",X"CE",X"BF",
		X"60",X"EE",X"C4",X"2A",X"0A",X"A6",X"52",X"26",X"F8",X"6A",X"53",X"26",X"F4",X"20",X"22",X"10",
		X"CE",X"BF",X"60",X"CC",X"E3",X"2F",X"DD",X"73",X"DE",X"5D",X"2B",X"03",X"CE",X"90",X"02",X"96",
		X"13",X"26",X"21",X"EE",X"C4",X"2A",X"1B",X"A6",X"52",X"27",X"F8",X"6A",X"53",X"26",X"F4",X"DF",
		X"5D",X"DF",X"21",X"6E",X"D8",X"F4",X"AE",X"E1",X"DE",X"21",X"AF",X"54",X"A7",X"53",X"6E",X"9F",
		X"90",X"73",X"DF",X"5D",X"96",X"13",X"27",X"FC",X"7E",X"E1",X"A4",X"34",X"17",X"1A",X"F0",X"8E",
		X"90",X"16",X"8D",X"08",X"8D",X"06",X"8D",X"04",X"8D",X"02",X"35",X"97",X"EC",X"81",X"2A",X"08",
		X"CC",X"B8",X"AB",X"ED",X"1E",X"7F",X"B8",X"AB",X"39",X"FE",X"B8",X"27",X"2A",X"33",X"E6",X"44",
		X"27",X"24",X"A1",X"43",X"25",X"2B",X"34",X"06",X"BE",X"03",X"22",X"EC",X"42",X"A3",X"84",X"ED",
		X"24",X"EC",X"02",X"ED",X"22",X"EC",X"06",X"ED",X"26",X"EC",X"44",X"ED",X"A4",X"5D",X"26",X"02",
		X"6F",X"44",X"31",X"28",X"35",X"06",X"33",X"46",X"11",X"83",X"B7",X"FB",X"23",X"D0",X"CE",X"00",
		X"00",X"FF",X"B8",X"27",X"39",X"DE",X"21",X"BD",X"E4",X"A5",X"24",X"27",X"6F",X"5E",X"86",X"01",
		X"BD",X"E3",X"46",X"8E",X"90",X"0E",X"11",X"A3",X"16",X"27",X"06",X"AE",X"16",X"2B",X"F7",X"20",
		X"12",X"EC",X"56",X"ED",X"16",X"11",X"93",X"0C",X"26",X"02",X"DD",X"0C",X"11",X"93",X"0A",X"26",
		X"02",X"DD",X"0A",X"EC",X"C4",X"8E",X"90",X"02",X"11",X"A3",X"84",X"27",X"07",X"AE",X"84",X"2B",
		X"F7",X"7E",X"E3",X"4E",X"ED",X"84",X"11",X"93",X"5D",X"26",X"02",X"9F",X"5D",X"DC",X"00",X"ED",
		X"C4",X"DF",X"00",X"9F",X"21",X"1F",X"13",X"7E",X"E3",X"4E",X"20",X"49",X"4E",X"46",X"45",X"52",
		X"4E",X"4F",X"20",X"2D",X"20",X"28",X"43",X"29",X"31",X"39",X"38",X"34",X"20",X"57",X"49",X"4C",
		X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",
		X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",X"34",X"46",X"8E",X"90",X"02",X"20",X"18",X"E6",X"61",
		X"E4",X"51",X"E1",X"E4",X"26",X"0E",X"11",X"93",X"21",X"27",X"09",X"CC",X"E3",X"B5",X"ED",X"54",
		X"86",X"01",X"A7",X"53",X"1F",X"31",X"EE",X"84",X"2B",X"E4",X"35",X"C6",X"DE",X"21",X"34",X"56",
		X"1F",X"21",X"10",X"9E",X"00",X"2B",X"04",X"1A",X"01",X"35",X"D6",X"EC",X"A4",X"DD",X"00",X"EC",
		X"C4",X"ED",X"A4",X"10",X"AF",X"C4",X"86",X"01",X"A7",X"33",X"AF",X"34",X"EC",X"E4",X"A7",X"31",
		X"E7",X"32",X"6F",X"28",X"4F",X"5F",X"ED",X"36",X"1C",X"FE",X"35",X"D6",X"39",X"9E",X"04",X"AF",
		X"56",X"DF",X"04",X"86",X"FF",X"A7",X"44",X"A7",X"46",X"CC",X"E4",X"8C",X"ED",X"C8",X"5A",X"ED",
		X"C8",X"58",X"ED",X"58",X"39",X"34",X"16",X"8E",X"90",X"0E",X"20",X"07",X"11",X"A3",X"16",X"27",
		X"0A",X"AE",X"16",X"EC",X"16",X"2B",X"F5",X"1C",X"FE",X"35",X"96",X"1A",X"01",X"35",X"96",X"34",
		X"06",X"4F",X"5F",X"DD",X"04",X"35",X"86",X"A6",X"C8",X"16",X"AB",X"C8",X"17",X"A7",X"48",X"9E",
		X"91",X"2A",X"02",X"8D",X"1C",X"9E",X"93",X"2A",X"02",X"8D",X"16",X"9E",X"95",X"2A",X"2B",X"8D",
		X"10",X"9E",X"97",X"2A",X"25",X"8D",X"0A",X"9E",X"99",X"2A",X"1F",X"8D",X"04",X"9E",X"9B",X"2A",
		X"19",X"EC",X"C8",X"1C",X"A0",X"88",X"1A",X"2D",X"11",X"E0",X"88",X"1B",X"2D",X"0C",X"A6",X"09",
		X"AB",X"48",X"A7",X"48",X"24",X"04",X"86",X"FF",X"A7",X"48",X"39",X"A6",X"C8",X"1C",X"AB",X"C8",
		X"1D",X"A7",X"48",X"E6",X"C8",X"57",X"E7",X"49",X"9E",X"91",X"2A",X"02",X"8D",X"1C",X"9E",X"93",
		X"2A",X"02",X"8D",X"16",X"9E",X"95",X"2A",X"44",X"8D",X"10",X"9E",X"97",X"2A",X"3E",X"8D",X"0A",
		X"9E",X"99",X"2A",X"38",X"8D",X"04",X"9E",X"9B",X"2A",X"32",X"9C",X"21",X"27",X"2E",X"EC",X"C8",
		X"1C",X"A0",X"88",X"1A",X"2D",X"26",X"E0",X"88",X"1B",X"2D",X"21",X"EC",X"88",X"1C",X"A0",X"C8",
		X"1A",X"2D",X"05",X"E0",X"C8",X"1B",X"2C",X"14",X"4F",X"E6",X"88",X"57",X"EB",X"49",X"E7",X"49",
		X"A6",X"09",X"AB",X"48",X"A7",X"48",X"24",X"04",X"86",X"FF",X"A7",X"48",X"39",X"34",X"06",X"F6",
		X"BF",X"FF",X"7F",X"BF",X"FF",X"7F",X"C8",X"00",X"7F",X"CB",X"A0",X"B7",X"C8",X"80",X"86",X"FF",
		X"B7",X"CB",X"A0",X"F7",X"BF",X"FF",X"F7",X"C8",X"00",X"35",X"86",X"34",X"06",X"F6",X"BF",X"FF",
		X"86",X"06",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"A6",X"E4",X"B7",X"C8",X"80",X"F7",X"BF",X"FF",
		X"F7",X"C8",X"00",X"35",X"86",X"F6",X"BF",X"FF",X"34",X"16",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",
		X"EC",X"84",X"ED",X"62",X"35",X"06",X"F7",X"BF",X"FF",X"F7",X"C8",X"00",X"35",X"86",X"B6",X"C9",
		X"80",X"B6",X"BF",X"FF",X"34",X"02",X"86",X"14",X"B7",X"C9",X"00",X"B6",X"CB",X"E0",X"84",X"C0",
		X"27",X"03",X"7E",X"E6",X"97",X"0C",X"1F",X"0A",X"20",X"B6",X"CB",X"E0",X"81",X"08",X"22",X"14",
		X"86",X"03",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"AD",X"9F",X"90",X"6F",X"86",X"01",X"B7",X"BF",
		X"FF",X"B7",X"C8",X"00",X"96",X"52",X"27",X"02",X"0A",X"52",X"DC",X"59",X"DD",X"5A",X"DC",X"57",
		X"DD",X"58",X"DC",X"55",X"DD",X"56",X"DC",X"53",X"DD",X"54",X"B6",X"C9",X"80",X"97",X"53",X"85",
		X"40",X"27",X"04",X"C6",X"78",X"D7",X"52",X"D6",X"53",X"DA",X"54",X"DA",X"55",X"DA",X"56",X"DA",
		X"57",X"DA",X"58",X"DA",X"59",X"DA",X"5A",X"DA",X"5B",X"D4",X"50",X"D7",X"51",X"94",X"54",X"9A",
		X"51",X"D6",X"50",X"97",X"50",X"53",X"1F",X"98",X"D4",X"50",X"C4",X"06",X"9A",X"50",X"43",X"84",
		X"38",X"A7",X"E2",X"EA",X"E0",X"34",X"04",X"DA",X"4F",X"D7",X"4F",X"86",X"01",X"B7",X"BF",X"FF",
		X"B7",X"C8",X"00",X"E6",X"E4",X"27",X"29",X"64",X"E4",X"64",X"E4",X"24",X"03",X"BD",X"F0",X"03",
		X"64",X"E4",X"24",X"03",X"BD",X"00",X"18",X"96",X"52",X"26",X"15",X"64",X"E4",X"24",X"03",X"BD",
		X"00",X"3C",X"64",X"E4",X"24",X"03",X"BD",X"00",X"3F",X"64",X"E4",X"24",X"03",X"BD",X"00",X"42",
		X"35",X"04",X"96",X"68",X"2A",X"11",X"DC",X"6B",X"83",X"00",X"01",X"2E",X"08",X"C6",X"06",X"BD",
		X"00",X"1E",X"CC",X"0E",X"10",X"DD",X"6B",X"10",X"DF",X"10",X"96",X"13",X"26",X"29",X"96",X"12",
		X"2F",X"0D",X"B6",X"CB",X"E0",X"84",X"C0",X"81",X"40",X"26",X"1C",X"0A",X"12",X"2E",X"18",X"9E",
		X"0E",X"30",X"02",X"8C",X"90",X"1E",X"25",X"12",X"0C",X"13",X"8E",X"90",X"14",X"9F",X"0E",X"0F",
		X"14",X"96",X"28",X"27",X"02",X"97",X"12",X"7E",X"E7",X"02",X"EE",X"84",X"60",X"84",X"9F",X"0E",
		X"96",X"14",X"8B",X"40",X"97",X"14",X"7A",X"C9",X"81",X"86",X"06",X"B7",X"BF",X"FF",X"B7",X"C8",
		X"00",X"20",X"02",X"34",X"3F",X"10",X"CE",X"C8",X"88",X"37",X"3F",X"29",X"F6",X"86",X"90",X"1F",
		X"8B",X"10",X"DE",X"10",X"1A",X"F0",X"7C",X"C9",X"81",X"B6",X"CB",X"E0",X"84",X"C0",X"90",X"14",
		X"26",X"AD",X"35",X"02",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"3B",X"8E",X"80",X"E0",X"BF",X"C8",
		X"84",X"8E",X"D0",X"00",X"BF",X"C8",X"82",X"CC",X"09",X"20",X"FD",X"C8",X"86",X"86",X"00",X"B7",
		X"C8",X"80",X"39",X"10",X"8E",X"D0",X"00",X"34",X"01",X"1A",X"F0",X"C6",X"40",X"A6",X"80",X"A7",
		X"A0",X"5A",X"26",X"F9",X"C6",X"20",X"30",X"88",X"E0",X"10",X"8C",X"D1",X"20",X"26",X"EE",X"CC",
		X"E7",X"0B",X"DD",X"6F",X"35",X"81",X"34",X"04",X"DC",X"1F",X"53",X"C5",X"09",X"26",X"05",X"53",
		X"46",X"56",X"20",X"09",X"53",X"C5",X"09",X"26",X"02",X"27",X"F5",X"44",X"56",X"DD",X"1F",X"44",
		X"35",X"84",X"34",X"06",X"A6",X"80",X"2B",X"04",X"D6",X"68",X"2A",X"10",X"91",X"4C",X"25",X"0C",
		X"97",X"4C",X"86",X"01",X"97",X"4B",X"9F",X"4D",X"A6",X"84",X"97",X"B6",X"35",X"86",X"34",X"02",
		X"B6",X"E7",X"B6",X"B7",X"C9",X"82",X"4F",X"97",X"4C",X"97",X"4B",X"97",X"B6",X"97",X"4D",X"97",
		X"4E",X"35",X"82",X"34",X"26",X"0D",X"68",X"2A",X"0D",X"E6",X"02",X"58",X"10",X"8E",X"90",X"A7",
		X"31",X"A5",X"EC",X"84",X"ED",X"A4",X"35",X"A6",X"34",X"10",X"8E",X"90",X"A7",X"6F",X"80",X"8C",
		X"90",X"B5",X"25",X"F9",X"35",X"90",X"00",X"00",X"01",X"02",X"03",X"04",X"04",X"06",X"06",X"06",
		X"06",X"06",X"07",X"7A",X"7A",X"17",X"0C",X"1E",X"1F",X"20",X"21",X"28",X"2E",X"32",X"A3",X"40",
		X"41",X"42",X"50",X"0D",X"08",X"09",X"0A",X"8C",X"8C",X"8C",X"0B",X"3E",X"89",X"4A",X"47",X"45",
		X"A3",X"0B",X"6F",X"5C",X"5C",X"79",X"75",X"76",X"A6",X"A1",X"52",X"A0",X"A4",X"1D",X"A7",X"4B",
		X"26",X"AE",X"75",X"34",X"02",X"B6",X"C9",X"86",X"84",X"C0",X"27",X"22",X"F6",X"CC",X"07",X"C4",
		X"0F",X"C1",X"09",X"27",X"0A",X"D6",X"E1",X"27",X"15",X"C1",X"02",X"24",X"02",X"84",X"7F",X"C6",
		X"01",X"85",X"80",X"26",X"05",X"85",X"40",X"27",X"05",X"5F",X"1A",X"01",X"35",X"82",X"1C",X"FE",
		X"35",X"82",X"96",X"9D",X"81",X"54",X"24",X"45",X"8E",X"A3",X"82",X"9F",X"29",X"86",X"01",X"D6",
		X"68",X"2B",X"10",X"BD",X"E7",X"F3",X"24",X"0B",X"86",X"01",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",
		X"7E",X"11",X"3E",X"5F",X"CE",X"BC",X"CA",X"1F",X"32",X"8E",X"00",X"00",X"AF",X"A1",X"AF",X"A1",
		X"AF",X"A1",X"AF",X"A1",X"AF",X"A1",X"AF",X"A1",X"AF",X"A1",X"AF",X"A1",X"10",X"8C",X"BE",X"1A",
		X"25",X"EA",X"BD",X"E8",X"6E",X"BD",X"E9",X"48",X"4C",X"91",X"A4",X"23",X"C2",X"39",X"34",X"06",
		X"8E",X"B8",X"AB",X"E6",X"E4",X"58",X"3A",X"3A",X"E6",X"80",X"27",X"03",X"5F",X"8D",X"23",X"33",
		X"C8",X"54",X"E6",X"80",X"27",X"04",X"C6",X"01",X"8D",X"18",X"33",X"C8",X"54",X"E6",X"80",X"27",
		X"04",X"C6",X"02",X"8D",X"0D",X"33",X"C8",X"54",X"E6",X"80",X"27",X"04",X"C6",X"03",X"8D",X"02",
		X"35",X"86",X"34",X"16",X"8E",X"BE",X"5A",X"4F",X"5F",X"ED",X"81",X"ED",X"81",X"ED",X"81",X"ED",
		X"81",X"8C",X"BE",X"AF",X"25",X"F3",X"10",X"8E",X"BE",X"5B",X"E6",X"E4",X"6C",X"A5",X"AE",X"62",
		X"A6",X"82",X"E6",X"A6",X"10",X"26",X"00",X"7E",X"C6",X"02",X"D7",X"9E",X"E7",X"A6",X"5A",X"E7",
		X"C6",X"0F",X"9F",X"8E",X"BE",X"5C",X"D6",X"9D",X"3A",X"96",X"9E",X"0C",X"9E",X"B7",X"BE",X"5A",
		X"A1",X"82",X"26",X"FC",X"8C",X"BE",X"5A",X"23",X"57",X"34",X"16",X"1F",X"10",X"83",X"BE",X"5B",
		X"58",X"58",X"49",X"C3",X"B8",X"AB",X"1F",X"01",X"E6",X"80",X"27",X"0D",X"A6",X"A5",X"26",X"09",
		X"96",X"9E",X"A7",X"A5",X"0C",X"9F",X"4A",X"A7",X"C5",X"E6",X"80",X"27",X"0D",X"A6",X"A5",X"26",
		X"09",X"96",X"9E",X"A7",X"A5",X"0C",X"9F",X"4A",X"A7",X"C5",X"E6",X"80",X"27",X"0D",X"A6",X"A5",
		X"26",X"09",X"96",X"9E",X"A7",X"A5",X"0C",X"9F",X"4A",X"A7",X"C5",X"E6",X"80",X"27",X"0D",X"A6",
		X"A5",X"26",X"09",X"96",X"9E",X"A7",X"A5",X"0C",X"9F",X"4A",X"A7",X"C5",X"35",X"16",X"20",X"A0",
		X"96",X"9F",X"10",X"26",X"FF",X"8B",X"35",X"96",X"34",X"42",X"CE",X"BC",X"CB",X"9E",X"29",X"96",
		X"9D",X"97",X"9F",X"10",X"8E",X"90",X"A0",X"A6",X"C4",X"E6",X"C8",X"54",X"DD",X"A0",X"A6",X"C9",
		X"00",X"A8",X"E6",X"C9",X"00",X"FC",X"DD",X"A2",X"5F",X"86",X"03",X"58",X"58",X"6D",X"A6",X"26",
		X"04",X"63",X"A6",X"CA",X"03",X"4A",X"2A",X"F3",X"E7",X"84",X"5F",X"8D",X"2A",X"25",X"1C",X"C6",
		X"40",X"8D",X"24",X"25",X"16",X"C6",X"80",X"8D",X"1E",X"25",X"10",X"C6",X"03",X"6D",X"A0",X"2B",
		X"06",X"1F",X"98",X"AA",X"84",X"A7",X"84",X"58",X"58",X"26",X"F2",X"33",X"41",X"30",X"01",X"0A",
		X"9F",X"26",X"B0",X"9F",X"29",X"35",X"C2",X"D7",X"9E",X"C6",X"7F",X"D1",X"A0",X"25",X"02",X"D6",
		X"A0",X"D1",X"A1",X"25",X"02",X"D6",X"A1",X"D1",X"A2",X"25",X"02",X"D6",X"A2",X"D1",X"A3",X"25",
		X"02",X"D6",X"A3",X"C1",X"7F",X"27",X"1A",X"86",X"03",X"E1",X"A6",X"26",X"0A",X"D6",X"9E",X"EA",
		X"84",X"E7",X"84",X"E6",X"A6",X"63",X"A6",X"04",X"9E",X"04",X"9E",X"4A",X"2A",X"EB",X"1C",X"FE",
		X"39",X"1A",X"01",X"39",X"32",X"7B",X"34",X"17",X"B6",X"BF",X"FF",X"A7",X"69",X"AE",X"6A",X"EC",
		X"81",X"ED",X"65",X"A6",X"80",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"AF",X"6A",X"CC",X"EA",X"04",
		X"ED",X"67",X"35",X"97",X"34",X"07",X"A6",X"63",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"35",X"07",
		X"32",X"61",X"39",X"96",X"71",X"26",X"04",X"AD",X"9F",X"E0",X"86",X"0A",X"71",X"2E",X"2F",X"86",
		X"07",X"97",X"71",X"96",X"72",X"0C",X"72",X"40",X"2E",X"3D",X"5F",X"8D",X"22",X"5C",X"D1",X"72",
		X"2D",X"F9",X"8D",X"1B",X"4C",X"91",X"72",X"2D",X"F9",X"8D",X"14",X"5A",X"2A",X"FB",X"FC",X"B8",
		X"18",X"C4",X"0F",X"DB",X"72",X"C1",X"10",X"25",X"05",X"FC",X"E0",X"86",X"DD",X"6F",X"39",X"34",
		X"06",X"BE",X"B8",X"18",X"48",X"48",X"48",X"30",X"86",X"30",X"86",X"30",X"85",X"31",X"89",X"04",
		X"00",X"A6",X"84",X"A7",X"A4",X"35",X"86",X"C6",X"03",X"3D",X"10",X"8E",X"EA",X"84",X"31",X"A5",
		X"A6",X"A4",X"97",X"71",X"BE",X"B8",X"18",X"30",X"89",X"04",X"00",X"EC",X"21",X"ED",X"84",X"88",
		X"80",X"C8",X"80",X"ED",X"88",X"10",X"39",X"10",X"1D",X"1E",X"04",X"1B",X"1C",X"1E",X"19",X"1A",
		X"34",X"46",X"F6",X"BF",X"FF",X"E7",X"E4",X"C6",X"05",X"F7",X"BF",X"FF",X"F7",X"C8",X"00",X"E6",
		X"61",X"CE",X"30",X"00",X"58",X"AB",X"D5",X"35",X"04",X"F7",X"BF",X"FF",X"F7",X"C8",X"00",X"35",
		X"C4",X"B6",X"BF",X"FF",X"34",X"02",X"86",X"05",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"C4",X"0F",
		X"58",X"AE",X"85",X"EC",X"81",X"1A",X"F0",X"10",X"BF",X"C8",X"84",X"31",X"A9",X"02",X"00",X"FD",
		X"C8",X"86",X"BF",X"C8",X"82",X"CC",X"12",X"00",X"F7",X"C8",X"81",X"B7",X"C8",X"80",X"1F",X"30",
		X"F7",X"C8",X"81",X"B7",X"C8",X"80",X"1C",X"EF",X"35",X"04",X"F7",X"BF",X"FF",X"F7",X"C8",X"00",
		X"39",X"F6",X"BF",X"FF",X"86",X"80",X"34",X"06",X"C6",X"06",X"F7",X"BF",X"FF",X"F7",X"C8",X"00",
		X"5F",X"1F",X"01",X"AB",X"82",X"5A",X"26",X"FB",X"6A",X"E4",X"26",X"F7",X"B0",X"EB",X"29",X"27",
		X"0F",X"10",X"9E",X"00",X"2A",X"0A",X"AE",X"A4",X"2A",X"04",X"1F",X"12",X"20",X"F8",X"6A",X"A4",
		X"35",X"06",X"F7",X"BF",X"FF",X"F7",X"C8",X"00",X"39",X"1F",X"00",X"00",X"FF",X"DF",X"75",X"CE",
		X"85",X"AE",X"A2",X"6F",X"AE",X"D1",X"BB",X"DA",X"EE",X"C1",X"00",X"00",X"0E",X"D1",X"0F",X"70",
		X"C0",X"D0",X"D8",X"89",X"E2",X"50",X"6A",X"DA",X"19",X"CC",X"00",X"00",X"AA",X"AB",X"CD",X"9B",
		X"BC",X"7A",X"AA",X"AB",X"CD",X"9B",X"BC",X"7A",X"CF",X"39",X"CF",X"59",X"CF",X"49",X"DF",X"2E",
		X"CC",X"7C",X"CC",X"BC",X"CC",X"AC",X"CC",X"9C",X"CC",X"8C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6F",X"4D",X"67",X"A4",X"69",X"BC",X"6F",X"EB",
		X"6B",X"32",X"6B",X"E3",X"6E",X"65",X"6A",X"8F",X"6D",X"B7",X"6C",X"21",X"6C",X"65",X"66",X"92",
		X"66",X"90",X"64",X"84",X"66",X"0F",X"66",X"65",X"68",X"BB",X"7E",X"60",X"E4",X"7E",X"63",X"6B",
		X"7E",X"60",X"00",X"7E",X"60",X"15",X"6D",X"48",X"6E",X"DB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E5",X"BE",X"E0",X"00",X"E0",X"00",X"E0",X"00",
		X"7E",X"F0",X"71",X"7E",X"F4",X"DF",X"7E",X"F6",X"3B",X"BD",X"BE",X"6F",X"49",X"00",X"05",X"39",
		X"BD",X"BE",X"6F",X"49",X"03",X"05",X"39",X"BD",X"BE",X"6F",X"49",X"06",X"05",X"39",X"BD",X"BE",
		X"6F",X"49",X"09",X"05",X"39",X"BD",X"BE",X"6F",X"49",X"0C",X"05",X"39",X"BD",X"BE",X"6F",X"49",
		X"0F",X"05",X"39",X"BD",X"BE",X"6F",X"49",X"12",X"05",X"39",X"BD",X"BE",X"6F",X"49",X"15",X"05",
		X"39",X"BD",X"BE",X"6F",X"49",X"18",X"05",X"39",X"BD",X"BE",X"6F",X"49",X"1B",X"05",X"39",X"BD",
		X"BE",X"6F",X"49",X"1E",X"05",X"39",X"BD",X"BE",X"6F",X"49",X"21",X"05",X"39",X"7E",X"BE",X"4E",
		X"7E",X"BE",X"10",X"7E",X"FA",X"23",X"7E",X"FF",X"6C",X"7E",X"F5",X"CE",X"7E",X"FA",X"13",X"F4",
		X"03",X"1A",X"FF",X"7F",X"CB",X"80",X"7F",X"CB",X"00",X"7F",X"CB",X"20",X"7F",X"C9",X"81",X"CC",
		X"00",X"3C",X"FD",X"C9",X"80",X"43",X"B7",X"C9",X"8C",X"86",X"02",X"20",X"2E",X"10",X"CE",X"BE",
		X"00",X"86",X"90",X"1F",X"8B",X"BD",X"F3",X"35",X"BD",X"F5",X"C7",X"25",X"15",X"BD",X"00",X"21",
		X"CC",X"01",X"99",X"8E",X"30",X"70",X"BD",X"E0",X"10",X"CC",X"02",X"99",X"8E",X"3A",X"90",X"BD",
		X"E0",X"10",X"10",X"8E",X"00",X"03",X"86",X"07",X"7E",X"F2",X"77",X"1A",X"3F",X"1F",X"8B",X"CE",
		X"00",X"00",X"8E",X"00",X"00",X"10",X"CE",X"BF",X"00",X"7F",X"C8",X"00",X"1F",X"30",X"53",X"C5",
		X"09",X"26",X"05",X"53",X"46",X"56",X"20",X"0B",X"53",X"C5",X"09",X"26",X"04",X"46",X"56",X"20",
		X"02",X"44",X"56",X"ED",X"81",X"1E",X"10",X"5D",X"26",X"16",X"C6",X"14",X"F7",X"C9",X"00",X"1F",
		X"B9",X"C1",X"FF",X"26",X"0A",X"F6",X"C9",X"80",X"C5",X"02",X"27",X"03",X"7E",X"F5",X"5A",X"5F",
		X"1E",X"10",X"11",X"8C",X"BF",X"03",X"26",X"07",X"8C",X"88",X"00",X"26",X"C1",X"20",X"1B",X"8C",
		X"C8",X"00",X"26",X"03",X"8E",X"D0",X"00",X"8C",X"E0",X"00",X"26",X"B2",X"8E",X"80",X"00",X"1E",
		X"04",X"C6",X"03",X"F7",X"C8",X"00",X"1E",X"04",X"20",X"A4",X"1F",X"32",X"8E",X"00",X"00",X"10",
		X"CE",X"BF",X"00",X"7F",X"C8",X"00",X"1F",X"20",X"53",X"C5",X"09",X"26",X"05",X"53",X"46",X"56",
		X"20",X"0B",X"53",X"C5",X"09",X"26",X"04",X"46",X"56",X"20",X"02",X"44",X"56",X"1F",X"02",X"A8",
		X"81",X"26",X"60",X"E8",X"1F",X"26",X"5C",X"1F",X"10",X"5D",X"26",X"15",X"C6",X"14",X"F7",X"C9",
		X"00",X"1F",X"B9",X"C1",X"FF",X"26",X"0A",X"F6",X"C9",X"80",X"C5",X"02",X"27",X"03",X"7E",X"F5",
		X"5A",X"11",X"8C",X"BF",X"03",X"26",X"07",X"8C",X"88",X"00",X"26",X"BA",X"20",X"1B",X"8C",X"C8",
		X"00",X"26",X"03",X"8E",X"D0",X"00",X"8C",X"E0",X"00",X"26",X"AB",X"8E",X"80",X"00",X"1E",X"04",
		X"C6",X"03",X"F7",X"C8",X"00",X"1E",X"04",X"20",X"9D",X"1F",X"23",X"1F",X"B8",X"81",X"FF",X"26",
		X"03",X"7E",X"F0",X"C2",X"4A",X"1F",X"8B",X"81",X"80",X"10",X"27",X"04",X"A7",X"4D",X"26",X"F1",
		X"7E",X"F0",X"8D",X"30",X"1E",X"11",X"8C",X"BF",X"03",X"27",X"1B",X"8C",X"CF",X"FF",X"22",X"0A",
		X"8C",X"C0",X"00",X"25",X"27",X"CE",X"04",X"40",X"20",X"56",X"CE",X"06",X"54",X"8C",X"D8",X"00",
		X"25",X"4E",X"33",X"41",X"20",X"4A",X"CE",X"05",X"78",X"85",X"F0",X"26",X"43",X"33",X"5F",X"4D",
		X"26",X"3E",X"33",X"5F",X"C5",X"F0",X"26",X"38",X"33",X"5F",X"20",X"34",X"4D",X"26",X"02",X"1F",
		X"98",X"1E",X"01",X"C6",X"14",X"F7",X"C9",X"00",X"80",X"03",X"24",X"F9",X"8B",X"03",X"1F",X"89",
		X"4F",X"58",X"58",X"58",X"1E",X"10",X"C6",X"FF",X"5C",X"48",X"24",X"FC",X"C8",X"03",X"3A",X"1F",
		X"10",X"8B",X"01",X"19",X"5A",X"2A",X"FA",X"8B",X"97",X"19",X"1F",X"89",X"86",X"01",X"1F",X"03",
		X"86",X"01",X"B7",X"C8",X"00",X"1F",X"30",X"10",X"CE",X"F2",X"2D",X"20",X"5E",X"1F",X"A8",X"10",
		X"CE",X"BE",X"00",X"11",X"83",X"01",X"99",X"22",X"04",X"10",X"CE",X"DF",X"FF",X"BD",X"F4",X"C9",
		X"C6",X"22",X"85",X"40",X"27",X"08",X"86",X"01",X"8E",X"30",X"70",X"BD",X"E0",X"10",X"86",X"03",
		X"8E",X"40",X"90",X"BD",X"E0",X"10",X"1F",X"30",X"8A",X"F0",X"C6",X"BB",X"BD",X"E0",X"17",X"1F",
		X"30",X"1F",X"98",X"C6",X"BB",X"BD",X"E0",X"17",X"1F",X"A8",X"85",X"40",X"26",X"03",X"7E",X"F5",
		X"77",X"10",X"8E",X"00",X"03",X"86",X"20",X"8E",X"58",X"00",X"30",X"1F",X"C6",X"14",X"F7",X"C9",
		X"00",X"8C",X"00",X"00",X"26",X"F4",X"4A",X"26",X"EE",X"6E",X"A4",X"1F",X"03",X"86",X"02",X"1F",
		X"8B",X"1F",X"30",X"10",X"8E",X"F2",X"9A",X"7E",X"F3",X"06",X"84",X"7F",X"B7",X"C9",X"8C",X"86",
		X"02",X"10",X"8E",X"F2",X"A7",X"20",X"D0",X"86",X"FF",X"B7",X"C9",X"8C",X"86",X"01",X"10",X"8E",
		X"F2",X"B4",X"20",X"C3",X"1F",X"30",X"1F",X"98",X"44",X"44",X"44",X"44",X"10",X"8E",X"F2",X"C2",
		X"20",X"44",X"86",X"02",X"10",X"8E",X"F2",X"CA",X"20",X"AD",X"86",X"FF",X"B7",X"C9",X"8C",X"86",
		X"01",X"10",X"8E",X"F2",X"D7",X"20",X"A0",X"1F",X"30",X"1F",X"98",X"10",X"8E",X"F2",X"E1",X"20",
		X"25",X"86",X"02",X"10",X"8E",X"F2",X"E9",X"20",X"8E",X"86",X"FF",X"B7",X"C9",X"8C",X"86",X"05",
		X"10",X"8E",X"F2",X"F6",X"20",X"81",X"1F",X"B8",X"4A",X"1F",X"8B",X"26",X"94",X"86",X"FF",X"B7",
		X"C9",X"8C",X"1F",X"30",X"6E",X"E4",X"84",X"0F",X"8E",X"F3",X"12",X"A6",X"86",X"B7",X"C9",X"8C",
		X"6E",X"A4",X"C0",X"F9",X"A4",X"B0",X"99",X"92",X"82",X"F8",X"80",X"90",X"88",X"83",X"C6",X"A1",
		X"86",X"8E",X"34",X"7F",X"10",X"FF",X"90",X"E6",X"10",X"CE",X"F3",X"2F",X"7E",X"F2",X"8B",X"10",
		X"FE",X"90",X"E6",X"35",X"FF",X"1A",X"3F",X"BD",X"F5",X"CE",X"4F",X"1F",X"8B",X"8E",X"F4",X"03",
		X"BD",X"FF",X"AB",X"EC",X"81",X"81",X"BF",X"27",X"F7",X"FD",X"C8",X"86",X"EC",X"84",X"FD",X"C8",
		X"84",X"E6",X"02",X"F7",X"C8",X"81",X"86",X"12",X"B7",X"C8",X"80",X"30",X"07",X"8C",X"F4",X"C8",
		X"25",X"DE",X"8E",X"F4",X"03",X"EC",X"81",X"81",X"BF",X"26",X"08",X"F7",X"BF",X"FF",X"F7",X"C8",
		X"00",X"20",X"F2",X"A6",X"06",X"81",X"00",X"27",X"46",X"A6",X"03",X"5F",X"1F",X"03",X"4F",X"EB",
		X"C0",X"4A",X"26",X"FB",X"BD",X"FA",X"13",X"25",X"3D",X"1E",X"03",X"A1",X"04",X"1E",X"03",X"26",
		X"ED",X"EE",X"1E",X"FF",X"C8",X"86",X"EE",X"84",X"FF",X"C8",X"84",X"E1",X"06",X"27",X"17",X"CC",
		X"12",X"22",X"F7",X"C8",X"81",X"B7",X"C8",X"80",X"1F",X"B8",X"4C",X"1F",X"8B",X"86",X"02",X"E6",
		X"05",X"BD",X"F3",X"22",X"20",X"09",X"CC",X"12",X"AA",X"F7",X"C8",X"81",X"B7",X"C8",X"80",X"30",
		X"07",X"8C",X"F4",X"C8",X"25",X"9F",X"86",X"01",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"1F",X"B8",
		X"4D",X"26",X"06",X"BD",X"FA",X"13",X"25",X"FB",X"39",X"1F",X"A8",X"43",X"85",X"C0",X"26",X"09",
		X"CC",X"01",X"22",X"8E",X"30",X"42",X"BD",X"E0",X"10",X"CC",X"04",X"22",X"8E",X"40",X"52",X"BD",
		X"E0",X"10",X"10",X"8E",X"F3",X"FB",X"86",X"07",X"7E",X"F2",X"77",X"BD",X"FA",X"13",X"25",X"FB",
		X"1A",X"01",X"39",X"90",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"80",X"10",X"40",
		X"99",X"00",X"00",X"00",X"00",X"18",X"06",X"38",X"C0",X"11",X"00",X"00",X"00",X"00",X"BF",X"05",
		X"0B",X"07",X"5C",X"AA",X"66",X"00",X"20",X"17",X"06",X"0B",X"07",X"5C",X"94",X"66",X"20",X"40",
		X"15",X"A4",X"0B",X"07",X"50",X"AA",X"66",X"40",X"60",X"13",X"30",X"0B",X"07",X"50",X"94",X"66",
		X"60",X"80",X"11",X"AF",X"BF",X"06",X"0B",X"07",X"74",X"AA",X"66",X"00",X"20",X"25",X"0C",X"0B",
		X"07",X"74",X"94",X"66",X"20",X"40",X"23",X"7E",X"0B",X"07",X"68",X"AA",X"66",X"40",X"60",X"21",
		X"44",X"0B",X"07",X"68",X"94",X"66",X"60",X"80",X"19",X"D1",X"BF",X"02",X"0B",X"07",X"74",X"B5",
		X"66",X"00",X"20",X"26",X"00",X"0B",X"07",X"74",X"9F",X"66",X"20",X"40",X"24",X"00",X"0B",X"07",
		X"68",X"B5",X"66",X"40",X"60",X"22",X"00",X"0B",X"07",X"68",X"9F",X"66",X"60",X"80",X"20",X"00",
		X"BF",X"01",X"0B",X"07",X"5C",X"B5",X"66",X"00",X"20",X"18",X"98",X"0B",X"07",X"5C",X"9F",X"66",
		X"20",X"40",X"16",X"E5",X"0B",X"07",X"50",X"B5",X"66",X"40",X"60",X"14",X"86",X"0B",X"07",X"50",
		X"9F",X"66",X"60",X"80",X"12",X"49",X"0B",X"07",X"3A",X"70",X"66",X"E0",X"F0",X"09",X"34",X"0B",
		X"07",X"3A",X"7B",X"66",X"F0",X"00",X"10",X"80",X"80",X"34",X"04",X"C6",X"90",X"1F",X"9B",X"C6",
		X"01",X"F7",X"BF",X"FF",X"F7",X"C8",X"00",X"BD",X"00",X"21",X"BD",X"F5",X"CE",X"35",X"84",X"10",
		X"CE",X"BE",X"00",X"86",X"90",X"1F",X"8B",X"86",X"01",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"4F",
		X"B7",X"CB",X"80",X"B7",X"C9",X"85",X"B7",X"C9",X"87",X"B7",X"C9",X"81",X"B7",X"C9",X"83",X"C6",
		X"04",X"FD",X"C9",X"84",X"FD",X"C9",X"86",X"FD",X"C9",X"80",X"C6",X"2C",X"43",X"FD",X"C9",X"82",
		X"B7",X"C9",X"82",X"BD",X"F5",X"CE",X"BD",X"00",X"21",X"B6",X"C9",X"80",X"46",X"10",X"25",X"05",
		X"10",X"1A",X"BF",X"1C",X"BF",X"86",X"FF",X"B7",X"C9",X"8C",X"BD",X"FF",X"AB",X"B6",X"C9",X"80",
		X"85",X"02",X"26",X"F6",X"BD",X"F3",X"35",X"86",X"00",X"BD",X"E0",X"33",X"C6",X"03",X"8E",X"70",
		X"00",X"BD",X"FF",X"AB",X"B6",X"C9",X"80",X"85",X"02",X"26",X"0F",X"30",X"1F",X"8C",X"00",X"00",
		X"26",X"EF",X"5A",X"26",X"E9",X"86",X"FF",X"7E",X"F0",X"BB",X"10",X"CE",X"BE",X"00",X"BD",X"F4",
		X"C9",X"86",X"01",X"BD",X"E0",X"33",X"8E",X"1A",X"0A",X"BD",X"FF",X"AB",X"B6",X"C9",X"80",X"85",
		X"02",X"26",X"F6",X"30",X"1F",X"26",X"F2",X"BD",X"F9",X"EB",X"CC",X"A5",X"5A",X"DD",X"C9",X"8D",
		X"46",X"BD",X"FF",X"0F",X"86",X"02",X"24",X"15",X"CC",X"03",X"59",X"8C",X"CD",X"00",X"22",X"01",
		X"5F",X"BD",X"F3",X"22",X"8D",X"31",X"86",X"03",X"5D",X"26",X"02",X"86",X"04",X"BD",X"00",X"21",
		X"BD",X"E0",X"33",X"BD",X"F9",X"EB",X"0F",X"C7",X"BD",X"FE",X"B3",X"BD",X"FE",X"BC",X"BD",X"FA",
		X"13",X"24",X"F8",X"4F",X"BD",X"FA",X"23",X"4F",X"BD",X"FF",X"0B",X"BD",X"F9",X"EB",X"BD",X"F8",
		X"EB",X"BD",X"F9",X"EB",X"7E",X"F6",X"8F",X"B6",X"F3",X"12",X"B7",X"C9",X"8C",X"39",X"34",X"56",
		X"8E",X"03",X"A7",X"B6",X"CB",X"E0",X"81",X"F9",X"27",X"04",X"30",X"1F",X"26",X"F5",X"CE",X"80",
		X"00",X"86",X"03",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"4F",X"5F",X"ED",X"C1",X"ED",X"C1",X"11",
		X"83",X"88",X"00",X"25",X"F6",X"CE",X"86",X"20",X"8E",X"F6",X"1B",X"EC",X"81",X"ED",X"C1",X"8C",
		X"F6",X"3B",X"25",X"F7",X"86",X"01",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"86",X"38",X"B7",X"CB",
		X"20",X"86",X"31",X"B7",X"CB",X"00",X"BD",X"FF",X"AB",X"35",X"D6",X"00",X"00",X"FB",X"AF",X"0F",
		X"A0",X"B0",X"A0",X"BF",X"A0",X"00",X"00",X"88",X"A8",X"4B",X"A0",X"0F",X"AF",X"FF",X"AF",X"F0",
		X"A0",X"4F",X"A0",X"38",X"AC",X"03",X"A8",X"03",X"A8",X"BF",X"A0",X"86",X"3C",X"B7",X"C9",X"81",
		X"B7",X"C9",X"85",X"B7",X"C9",X"87",X"86",X"2C",X"B7",X"C9",X"83",X"86",X"3F",X"1F",X"8A",X"86",
		X"8F",X"7E",X"F0",X"BB",X"10",X"CE",X"BE",X"00",X"86",X"90",X"1F",X"8B",X"BD",X"F3",X"35",X"25",
		X"1B",X"86",X"90",X"1F",X"8B",X"BD",X"FF",X"0F",X"24",X"17",X"86",X"04",X"8C",X"CD",X"00",X"23",
		X"02",X"86",X"03",X"BD",X"00",X"21",X"BD",X"F5",X"CE",X"BD",X"E0",X"33",X"BD",X"FF",X"AB",X"20",
		X"FB",X"BD",X"00",X"21",X"8D",X"5F",X"10",X"8E",X"F6",X"3B",X"86",X"04",X"7E",X"F2",X"77",X"BD",
		X"00",X"60",X"BD",X"F9",X"EB",X"BD",X"F7",X"4B",X"BD",X"F9",X"EB",X"CC",X"0F",X"D0",X"8D",X"12",
		X"CC",X"F0",X"D0",X"8D",X"0D",X"CC",X"00",X"DF",X"8D",X"08",X"8D",X"39",X"BD",X"F9",X"EB",X"7E",
		X"FA",X"31",X"1F",X"01",X"86",X"03",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"BF",X"86",X"22",X"86",
		X"01",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"8E",X"11",X"11",X"1F",X"12",X"1F",X"10",X"CE",X"90",
		X"00",X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"BD",X"FF",X"AB",X"11",X"83",X"90",X"00",
		X"25",X"EF",X"7E",X"F9",X"EB",X"86",X"03",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"8E",X"86",X"20",
		X"10",X"8E",X"F7",X"2B",X"EC",X"A1",X"ED",X"81",X"BD",X"FF",X"AB",X"8C",X"86",X"60",X"25",X"F4",
		X"86",X"01",X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"4F",X"5F",X"1F",X"01",X"9F",X"C5",X"30",X"89",
		X"0F",X"00",X"ED",X"83",X"BD",X"FF",X"AB",X"9C",X"C5",X"26",X"F7",X"30",X"89",X"08",X"00",X"4D",
		X"26",X"03",X"8E",X"0D",X"00",X"C3",X"11",X"11",X"24",X"E2",X"39",X"00",X"00",X"00",X"00",X"FF",
		X"DF",X"FF",X"DF",X"0F",X"D0",X"0F",X"D0",X"F0",X"D0",X"F0",X"D0",X"00",X"DF",X"00",X"DF",X"FF",
		X"D0",X"FF",X"D0",X"F0",X"DF",X"F0",X"DF",X"0F",X"DF",X"0F",X"DF",X"BD",X"00",X"21",X"86",X"03",
		X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"CC",X"FF",X"DF",X"FD",X"86",X"22",X"CC",X"00",X"DF",X"FD",
		X"86",X"24",X"CC",X"F0",X"D0",X"FD",X"86",X"26",X"CC",X"0F",X"D0",X"FD",X"86",X"28",X"7F",X"BF",
		X"FF",X"7F",X"C8",X"00",X"10",X"8E",X"F8",X"6B",X"86",X"01",X"AE",X"A4",X"BD",X"FF",X"AB",X"A7",
		X"80",X"AC",X"22",X"26",X"FA",X"31",X"24",X"10",X"8C",X"F8",X"93",X"26",X"ED",X"86",X"11",X"10",
		X"8E",X"F8",X"4B",X"AE",X"A4",X"9F",X"C5",X"A7",X"84",X"0C",X"C5",X"BD",X"FF",X"AB",X"9E",X"C5",
		X"AC",X"22",X"26",X"F3",X"31",X"24",X"10",X"8C",X"F8",X"6B",X"26",X"E7",X"10",X"8E",X"F8",X"93",
		X"AE",X"A4",X"9F",X"C5",X"A6",X"24",X"A7",X"84",X"0C",X"C5",X"BD",X"FF",X"AB",X"9E",X"C5",X"AC",
		X"22",X"26",X"F3",X"31",X"25",X"10",X"8C",X"F8",X"CF",X"26",X"E5",X"10",X"8E",X"F8",X"CF",X"AE",
		X"A4",X"A6",X"24",X"A7",X"80",X"BD",X"FF",X"AB",X"AC",X"22",X"26",X"F7",X"31",X"25",X"10",X"8C",
		X"F8",X"E3",X"26",X"EB",X"86",X"21",X"B7",X"3F",X"7F",X"86",X"20",X"B7",X"8C",X"7F",X"8E",X"47",
		X"0D",X"A6",X"84",X"84",X"F0",X"8A",X"02",X"BD",X"FF",X"AB",X"A7",X"80",X"8C",X"47",X"6D",X"26",
		X"F0",X"8E",X"47",X"90",X"A6",X"84",X"84",X"F0",X"8A",X"02",X"BD",X"FF",X"AB",X"A7",X"80",X"8C",
		X"47",X"F3",X"26",X"F0",X"8E",X"0A",X"19",X"10",X"8E",X"F8",X"E3",X"9F",X"C5",X"9E",X"C5",X"A6",
		X"84",X"84",X"F0",X"8A",X"01",X"A7",X"84",X"D6",X"C6",X"CB",X"22",X"25",X"04",X"D7",X"C6",X"20",
		X"EC",X"C6",X"19",X"D7",X"C6",X"E6",X"A0",X"D7",X"C5",X"10",X"8C",X"F8",X"EC",X"26",X"DE",X"C6",
		X"01",X"F7",X"BF",X"FF",X"F7",X"C8",X"00",X"BD",X"FF",X"AB",X"39",X"05",X"09",X"8D",X"09",X"05",
		X"2A",X"8D",X"2A",X"05",X"4C",X"8D",X"4C",X"05",X"6E",X"8D",X"6E",X"05",X"90",X"8D",X"90",X"05",
		X"B4",X"8D",X"B4",X"05",X"D6",X"8D",X"D6",X"05",X"F6",X"8D",X"F6",X"05",X"09",X"05",X"F6",X"11",
		X"09",X"11",X"F6",X"20",X"09",X"20",X"F6",X"30",X"09",X"30",X"F6",X"3F",X"09",X"3F",X"F6",X"4F",
		X"09",X"4F",X"F6",X"5E",X"09",X"5E",X"F6",X"6E",X"09",X"6E",X"F6",X"7D",X"09",X"7D",X"F6",X"8C",
		X"09",X"8C",X"F6",X"42",X"07",X"4D",X"07",X"44",X"42",X"08",X"4D",X"08",X"44",X"42",X"09",X"4D",
		X"09",X"00",X"42",X"0A",X"4D",X"0A",X"33",X"42",X"0B",X"4D",X"0B",X"33",X"42",X"F4",X"4D",X"F4",
		X"33",X"42",X"F5",X"4D",X"F5",X"33",X"42",X"F6",X"4D",X"F6",X"00",X"42",X"F7",X"4D",X"F7",X"44",
		X"42",X"F8",X"4D",X"F8",X"44",X"05",X"7F",X"3F",X"7F",X"22",X"50",X"7F",X"8C",X"7F",X"22",X"04",
		X"70",X"04",X"8F",X"43",X"05",X"70",X"05",X"8F",X"00",X"8C",X"70",X"8C",X"8F",X"00",X"8D",X"70",
		X"8D",X"8F",X"34",X"18",X"28",X"37",X"47",X"56",X"66",X"76",X"85",X"86",X"0A",X"97",X"C5",X"BD",
		X"00",X"21",X"86",X"05",X"BD",X"E0",X"33",X"CE",X"90",X"E8",X"6F",X"C0",X"11",X"83",X"90",X"F1",
		X"23",X"F8",X"CE",X"F9",X"73",X"10",X"8E",X"90",X"E9",X"C6",X"2C",X"AE",X"C1",X"6F",X"84",X"4F",
		X"A7",X"1F",X"A6",X"C0",X"A7",X"84",X"AE",X"C1",X"A6",X"A4",X"34",X"02",X"A6",X"84",X"A8",X"C0",
		X"A7",X"A4",X"A8",X"E0",X"97",X"E8",X"A6",X"A0",X"1A",X"01",X"46",X"8D",X"13",X"44",X"26",X"FB",
		X"11",X"83",X"F9",X"EB",X"25",X"D5",X"BD",X"FA",X"13",X"24",X"C7",X"0A",X"C5",X"26",X"C3",X"39",
		X"34",X"36",X"BD",X"FF",X"AB",X"A6",X"41",X"27",X"24",X"A6",X"42",X"1F",X"01",X"86",X"BB",X"24",
		X"02",X"86",X"11",X"CB",X"07",X"E7",X"61",X"1F",X"89",X"A6",X"C4",X"BD",X"E0",X"25",X"A6",X"41",
		X"BD",X"E0",X"2C",X"96",X"E8",X"44",X"24",X"05",X"86",X"01",X"BD",X"FF",X"0B",X"33",X"43",X"04",
		X"E8",X"35",X"B6",X"C9",X"81",X"34",X"C9",X"80",X"00",X"0F",X"FF",X"43",X"10",X"FF",X"43",X"12",
		X"FF",X"3A",X"13",X"FF",X"41",X"14",X"FF",X"3F",X"11",X"FF",X"40",X"15",X"FF",X"3E",X"00",X"00",
		X"00",X"C9",X"85",X"34",X"C9",X"84",X"FF",X"18",X"F1",X"3C",X"19",X"F1",X"3D",X"1A",X"F1",X"3A",
		X"1B",X"F1",X"3B",X"1C",X"F1",X"3C",X"1D",X"F1",X"3D",X"5B",X"F1",X"39",X"5C",X"F1",X"3A",X"C9",
		X"87",X"34",X"C9",X"86",X"00",X"5D",X"F1",X"41",X"5D",X"F2",X"41",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"FF",X"3A",X"17",X"FF",X"3A",X"C9",X"85",X"3C",
		X"C9",X"84",X"FF",X"18",X"F2",X"3C",X"19",X"F2",X"3D",X"1A",X"F2",X"3A",X"1B",X"F2",X"3B",X"1C",
		X"F2",X"3C",X"1D",X"F2",X"3D",X"5B",X"F2",X"39",X"5C",X"F2",X"3A",X"86",X"01",X"B7",X"BF",X"FF",
		X"B7",X"C8",X"00",X"BD",X"FA",X"13",X"25",X"06",X"86",X"01",X"8D",X"27",X"20",X"ED",X"86",X"01",
		X"B7",X"BF",X"FF",X"B7",X"C8",X"00",X"BD",X"00",X"21",X"86",X"01",X"8D",X"16",X"BD",X"FA",X"13",
		X"25",X"F7",X"39",X"BD",X"FF",X"AB",X"B6",X"C9",X"80",X"85",X"02",X"27",X"03",X"1A",X"01",X"39",
		X"1C",X"FE",X"39",X"8E",X"01",X"00",X"BD",X"FF",X"AB",X"30",X"1F",X"26",X"F9",X"4A",X"2A",X"F3",
		X"39",X"86",X"90",X"1F",X"8B",X"BD",X"F5",X"CE",X"8D",X"C4",X"86",X"06",X"BD",X"E0",X"33",X"CE",
		X"CD",X"02",X"8E",X"1A",X"30",X"86",X"20",X"34",X"12",X"C6",X"88",X"BD",X"E0",X"10",X"1E",X"31",
		X"BD",X"00",X"27",X"C5",X"F0",X"26",X"08",X"CA",X"F0",X"C5",X"0F",X"26",X"02",X"CA",X"0F",X"1F",
		X"98",X"43",X"34",X"06",X"BD",X"00",X"2A",X"6D",X"E0",X"26",X"12",X"85",X"F0",X"26",X"0E",X"8A",
		X"F0",X"85",X"0F",X"26",X"08",X"8A",X"0F",X"C5",X"F0",X"26",X"02",X"CA",X"F0",X"1F",X"02",X"1E",
		X"31",X"1F",X"10",X"86",X"6A",X"1F",X"01",X"35",X"02",X"C6",X"88",X"BD",X"E0",X"17",X"BD",X"FF",
		X"AB",X"1F",X"20",X"34",X"04",X"C6",X"88",X"BD",X"E0",X"17",X"35",X"02",X"BD",X"E0",X"17",X"BD",
		X"FF",X"AB",X"35",X"12",X"30",X"0E",X"4C",X"11",X"83",X"CD",X"3E",X"23",X"9A",X"86",X"2B",X"C6",
		X"88",X"BD",X"E0",X"10",X"1F",X"10",X"86",X"6E",X"1F",X"01",X"1E",X"31",X"8E",X"CD",X"20",X"BD",
		X"00",X"27",X"D7",X"CE",X"BD",X"00",X"2A",X"DD",X"CF",X"8E",X"CD",X"3E",X"BD",X"00",X"27",X"D7",
		X"D1",X"BD",X"00",X"2A",X"DD",X"D2",X"1E",X"31",X"8D",X"29",X"C6",X"88",X"85",X"F0",X"26",X"02",
		X"8A",X"F0",X"BD",X"E0",X"17",X"34",X"10",X"30",X"1C",X"86",X"2E",X"BD",X"E0",X"09",X"35",X"10",
		X"86",X"2E",X"BD",X"E0",X"09",X"96",X"D0",X"BD",X"E0",X"17",X"BD",X"FF",X"AB",X"BD",X"F9",X"EB",
		X"7E",X"FC",X"E5",X"34",X"30",X"8D",X"66",X"DC",X"CE",X"27",X"0C",X"86",X"99",X"34",X"02",X"97",
		X"D0",X"0F",X"CF",X"0F",X"CE",X"20",X"3C",X"96",X"D0",X"34",X"02",X"DC",X"CB",X"DD",X"CE",X"96",
		X"CD",X"97",X"D0",X"4F",X"5F",X"DD",X"CB",X"97",X"CD",X"86",X"04",X"08",X"D0",X"09",X"CF",X"09",
		X"CE",X"09",X"CD",X"4A",X"26",X"F5",X"8E",X"90",X"D1",X"10",X"8E",X"90",X"D1",X"CE",X"90",X"D1",
		X"8D",X"13",X"DC",X"CD",X"DD",X"D4",X"DC",X"CF",X"DD",X"D6",X"8E",X"90",X"D8",X"8D",X"06",X"8D",
		X"04",X"8D",X"20",X"35",X"B2",X"34",X"70",X"C6",X"04",X"20",X"04",X"34",X"70",X"C6",X"03",X"1C",
		X"FE",X"A6",X"82",X"A9",X"A2",X"19",X"A7",X"C2",X"5A",X"26",X"F6",X"35",X"F0",X"4F",X"5F",X"DD",
		X"CB",X"97",X"CD",X"DC",X"D1",X"26",X"0B",X"96",X"D3",X"26",X"07",X"4F",X"5F",X"DD",X"CE",X"97",
		X"D0",X"39",X"86",X"07",X"97",X"D4",X"8E",X"90",X"CE",X"10",X"8E",X"90",X"D4",X"CE",X"90",X"D8",
		X"8D",X"29",X"0A",X"D4",X"26",X"02",X"20",X"23",X"86",X"04",X"08",X"D0",X"09",X"CF",X"09",X"CE",
		X"09",X"CD",X"09",X"CC",X"09",X"CB",X"4A",X"26",X"F1",X"8D",X"B0",X"25",X"02",X"20",X"E3",X"DC",
		X"D5",X"DD",X"CB",X"96",X"D7",X"97",X"CD",X"0C",X"D0",X"20",X"EE",X"34",X"20",X"C6",X"03",X"86",
		X"99",X"A0",X"A2",X"A7",X"A4",X"5A",X"26",X"F7",X"10",X"AE",X"E4",X"C6",X"03",X"1A",X"01",X"A6",
		X"3F",X"89",X"00",X"19",X"A7",X"A2",X"5A",X"26",X"F6",X"35",X"A0",X"2D",X"6A",X"1A",X"20",X"CC",
		X"00",X"FE",X"42",X"00",X"99",X"FD",X"FB",X"FE",X"00",X"2E",X"6A",X"1A",X"29",X"CC",X"02",X"FE",
		X"37",X"01",X"99",X"FD",X"FB",X"FD",X"FE",X"2F",X"6A",X"1A",X"32",X"CC",X"04",X"FE",X"29",X"00",
		X"01",X"FD",X"FB",X"FD",X"FE",X"30",X"6A",X"1A",X"3B",X"CC",X"06",X"FE",X"4E",X"00",X"09",X"FE",
		X"01",X"FD",X"FE",X"31",X"6A",X"22",X"44",X"CC",X"08",X"FE",X"37",X"00",X"99",X"FD",X"FB",X"FD",
		X"FE",X"32",X"6A",X"22",X"4D",X"CC",X"0A",X"FE",X"37",X"00",X"99",X"FD",X"FB",X"FD",X"FE",X"33",
		X"6A",X"22",X"56",X"CC",X"0C",X"FE",X"37",X"00",X"99",X"FD",X"FB",X"FD",X"FE",X"34",X"6A",X"22",
		X"5F",X"CC",X"0E",X"FE",X"37",X"01",X"99",X"FD",X"FB",X"FD",X"FE",X"35",X"6A",X"22",X"68",X"CC",
		X"10",X"FE",X"37",X"00",X"99",X"FD",X"FB",X"FD",X"FE",X"36",X"6A",X"22",X"71",X"CC",X"12",X"FE",
		X"37",X"00",X"99",X"FD",X"FB",X"FD",X"FE",X"37",X"6A",X"1A",X"7A",X"CC",X"14",X"FE",X"37",X"00",
		X"09",X"FD",X"FB",X"FE",X"0C",X"38",X"6A",X"1A",X"83",X"CC",X"16",X"FE",X"37",X"03",X"20",X"FD",
		X"FB",X"FD",X"FE",X"A6",X"6A",X"1A",X"8C",X"CC",X"18",X"FE",X"29",X"00",X"01",X"FD",X"FB",X"FD",
		X"FE",X"39",X"6A",X"1A",X"95",X"CC",X"1A",X"FE",X"29",X"00",X"01",X"FD",X"FB",X"FD",X"FE",X"3A",
		X"6A",X"1A",X"9E",X"CC",X"1C",X"FE",X"29",X"00",X"01",X"FD",X"FB",X"FD",X"FE",X"3B",X"6A",X"1A",
		X"A7",X"CC",X"1E",X"FE",X"29",X"00",X"01",X"FD",X"FB",X"FD",X"FE",X"3C",X"6A",X"1A",X"B0",X"CC",
		X"20",X"FE",X"29",X"00",X"01",X"FD",X"FB",X"FD",X"FE",X"3D",X"6A",X"1A",X"B9",X"CC",X"22",X"FE",
		X"29",X"00",X"01",X"FD",X"FB",X"FD",X"FE",X"3E",X"6A",X"1A",X"C2",X"CC",X"24",X"FE",X"29",X"00",
		X"01",X"FE",X"00",X"FD",X"FE",X"8E",X"CC",X"1A",X"6F",X"80",X"8C",X"CC",X"26",X"25",X"F9",X"BD",
		X"F9",X"FE",X"86",X"07",X"BD",X"E0",X"33",X"CE",X"FB",X"DB",X"5F",X"BD",X"FD",X"DA",X"33",X"4E",
		X"11",X"83",X"FC",X"E5",X"25",X"F4",X"86",X"08",X"BD",X"E0",X"3A",X"CE",X"FB",X"DB",X"86",X"0C",
		X"97",X"E8",X"97",X"E9",X"C6",X"33",X"BD",X"FD",X"DA",X"BD",X"FA",X"13",X"24",X"06",X"BD",X"F9",
		X"FE",X"7E",X"00",X"0C",X"D6",X"E8",X"2B",X"02",X"0A",X"E8",X"D6",X"E9",X"2B",X"02",X"0A",X"E9",
		X"86",X"01",X"BD",X"FA",X"23",X"BD",X"00",X"57",X"C5",X"0F",X"27",X"1E",X"96",X"E8",X"2E",X"D9",
		X"86",X"0A",X"97",X"E8",X"34",X"04",X"5F",X"BD",X"FD",X"DA",X"35",X"04",X"C5",X"03",X"27",X"05",
		X"AD",X"D8",X"0C",X"20",X"BF",X"AD",X"D8",X"0A",X"20",X"BA",X"0F",X"E8",X"C5",X"F0",X"26",X"05",
		X"0F",X"E9",X"7E",X"FD",X"19",X"96",X"E9",X"2E",X"F9",X"86",X"14",X"0D",X"E9",X"2B",X"02",X"86",
		X"03",X"97",X"E9",X"34",X"04",X"C6",X"33",X"AD",X"D8",X"06",X"86",X"01",X"BD",X"FA",X"23",X"AE",
		X"44",X"BD",X"00",X"24",X"35",X"04",X"C5",X"30",X"27",X"0D",X"A1",X"49",X"25",X"04",X"A6",X"49",
		X"20",X"10",X"8B",X"01",X"19",X"20",X"0B",X"A1",X"48",X"22",X"04",X"A6",X"48",X"20",X"03",X"8B",
		X"99",X"19",X"AE",X"44",X"BD",X"00",X"2D",X"C6",X"11",X"AD",X"D8",X"06",X"11",X"83",X"FC",X"05",
		X"26",X"B0",X"34",X"40",X"8D",X"0E",X"8D",X"0C",X"8D",X"0A",X"8D",X"08",X"8D",X"06",X"8D",X"04",
		X"35",X"40",X"20",X"9E",X"34",X"04",X"33",X"4E",X"5F",X"AD",X"D8",X"06",X"AE",X"44",X"A6",X"A0",
		X"BD",X"00",X"2D",X"C6",X"11",X"AD",X"D8",X"06",X"35",X"84",X"F7",X"C8",X"81",X"EC",X"42",X"4F",
		X"5A",X"FD",X"C8",X"84",X"CC",X"90",X"07",X"FD",X"C8",X"86",X"86",X"12",X"B7",X"C8",X"80",X"A6",
		X"C4",X"AE",X"42",X"C6",X"11",X"BD",X"E0",X"25",X"6E",X"D8",X"06",X"33",X"4E",X"39",X"33",X"52",
		X"39",X"B6",X"CC",X"07",X"84",X"0F",X"27",X"F3",X"CE",X"FC",X"67",X"39",X"B6",X"CC",X"07",X"84",
		X"0F",X"27",X"EB",X"CE",X"FC",X"05",X"39",X"BD",X"FF",X"AB",X"AE",X"44",X"BD",X"00",X"24",X"34",
		X"06",X"EC",X"42",X"A6",X"41",X"1F",X"01",X"35",X"86",X"8D",X"EC",X"4D",X"27",X"04",X"86",X"41",
		X"20",X"02",X"86",X"08",X"7E",X"E0",X"25",X"8D",X"DE",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"7E",
		X"E0",X"2C",X"8D",X"F3",X"86",X"2D",X"BD",X"E0",X"1E",X"86",X"30",X"7E",X"E0",X"1E",X"8D",X"E7",
		X"84",X"0F",X"34",X"02",X"10",X"8E",X"FE",X"6D",X"31",X"A6",X"48",X"31",X"A6",X"48",X"31",X"A6",
		X"A6",X"A0",X"27",X"07",X"30",X"89",X"04",X"00",X"BD",X"E0",X"25",X"35",X"82",X"5F",X"01",X"04",
		X"01",X"01",X"00",X"00",X"00",X"01",X"04",X"01",X"02",X"04",X"00",X"00",X"06",X"00",X"01",X"01",
		X"00",X"00",X"00",X"01",X"04",X"01",X"01",X"00",X"00",X"00",X"01",X"16",X"06",X"02",X"00",X"00",
		X"00",X"01",X"04",X"01",X"02",X"00",X"00",X"00",X"01",X"00",X"04",X"01",X"00",X"00",X"00",X"01",
		X"00",X"02",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"02",X"00",X"00",X"5A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"BD",X"00",X"21",X"CC",X"01",X"01",X"DD",X"E9",X"39",X"4F",X"8D",X"4C",X"86",
		X"09",X"BD",X"FA",X"23",X"DC",X"E9",X"8D",X"43",X"8E",X"3A",X"80",X"CC",X"1E",X"99",X"BD",X"E0",
		X"10",X"96",X"EA",X"8A",X"F0",X"34",X"10",X"BD",X"E0",X"17",X"35",X"20",X"86",X"40",X"97",X"E8",
		X"86",X"01",X"BD",X"FA",X"23",X"BD",X"FA",X"13",X"25",X"04",X"0A",X"E8",X"26",X"F2",X"96",X"C7",
		X"26",X"06",X"B6",X"C9",X"80",X"46",X"24",X"12",X"1F",X"21",X"96",X"EA",X"8A",X"F0",X"5F",X"BD",
		X"E0",X"17",X"DC",X"E9",X"5C",X"48",X"25",X"AE",X"DD",X"E9",X"39",X"B7",X"C9",X"82",X"39",X"8E",
		X"CC",X"00",X"10",X"8E",X"90",X"00",X"A6",X"80",X"A7",X"A0",X"8C",X"D0",X"00",X"26",X"F7",X"C6",
		X"06",X"DE",X"C9",X"10",X"9E",X"C8",X"8E",X"CC",X"00",X"BD",X"FF",X"6C",X"A7",X"80",X"8D",X"7B",
		X"8C",X"D0",X"00",X"26",X"F4",X"10",X"9F",X"C8",X"DF",X"C9",X"8E",X"CC",X"00",X"BD",X"FF",X"6C",
		X"A8",X"80",X"84",X"0F",X"26",X"21",X"8D",X"63",X"8C",X"D0",X"00",X"26",X"F0",X"5A",X"26",X"D1",
		X"8D",X"03",X"1C",X"FE",X"39",X"CE",X"90",X"00",X"10",X"8E",X"CC",X"00",X"A6",X"C0",X"A7",X"A0",
		X"10",X"8C",X"D0",X"00",X"26",X"F6",X"39",X"8D",X"EC",X"1A",X"01",X"39",X"34",X"04",X"D6",X"C8",
		X"86",X"03",X"3D",X"CB",X"11",X"96",X"CA",X"44",X"44",X"44",X"98",X"CA",X"44",X"06",X"C9",X"06",
		X"CA",X"DB",X"CA",X"D9",X"C9",X"D7",X"C8",X"96",X"C8",X"35",X"84",X"28",X"43",X"29",X"31",X"39",
		X"38",X"34",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",
		X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"6E",X"9F",X"EF",X"F8",X"34",X"03",X"86",X"14",X"B7",
		X"C9",X"00",X"35",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A7",X"F0",X"00",X"F0",X"00",X"F0",X"00");
		

begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
