library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity inferno_bank_c is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of inferno_bank_c is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3F",X"3F",X"3F",X"7E",X"02",X"77",X"7E",X"02",X"F4",X"7E",X"01",X"10",X"7E",X"01",X"99",X"7E",
		X"05",X"0E",X"7E",X"03",X"56",X"7E",X"03",X"36",X"7E",X"03",X"02",X"7E",X"06",X"5F",X"7E",X"06",
		X"59",X"7E",X"06",X"09",X"7E",X"06",X"2A",X"7E",X"06",X"3B",X"7E",X"06",X"39",X"7E",X"06",X"43",
		X"7E",X"06",X"51",X"7E",X"06",X"4F",X"7E",X"06",X"98",X"7E",X"08",X"20",X"7E",X"08",X"42",X"7E",
		X"08",X"3C",X"7E",X"08",X"36",X"7E",X"08",X"9F",X"7E",X"08",X"B5",X"7E",X"08",X"CA",X"7E",X"09",
		X"38",X"7E",X"0A",X"32",X"7E",X"0B",X"B1",X"7E",X"00",X"63",X"7E",X"00",X"6F",X"7E",X"00",X"5D",
		X"7E",X"0F",X"57",X"34",X"72",X"CE",X"90",X"F2",X"C6",X"34",X"B6",X"C9",X"86",X"20",X"0B",X"34",
		X"72",X"CE",X"90",X"F8",X"C6",X"3C",X"B6",X"C9",X"86",X"44",X"7D",X"C9",X"80",X"2A",X"01",X"4F",
		X"84",X"01",X"F7",X"C9",X"85",X"F6",X"C9",X"84",X"C8",X"FF",X"34",X"06",X"AA",X"42",X"EA",X"43",
		X"AA",X"44",X"EA",X"45",X"A4",X"C4",X"E4",X"41",X"ED",X"C4",X"EC",X"E4",X"A4",X"42",X"E4",X"43",
		X"A4",X"44",X"E4",X"45",X"AA",X"C4",X"EA",X"41",X"ED",X"C4",X"EC",X"42",X"ED",X"44",X"35",X"06",
		X"ED",X"42",X"E6",X"C4",X"58",X"58",X"58",X"58",X"C4",X"10",X"EA",X"41",X"35",X"F2",X"0D",X"E4",
		X"27",X"3E",X"BD",X"11",X"32",X"86",X"04",X"BD",X"E0",X"7D",X"BD",X"00",X"21",X"8E",X"20",X"20",
		X"86",X"55",X"C6",X"11",X"BD",X"E0",X"10",X"8E",X"14",X"CA",X"86",X"57",X"C6",X"99",X"BD",X"E0",
		X"25",X"BE",X"11",X"09",X"BD",X"E0",X"75",X"6F",X"C8",X"30",X"86",X"1E",X"BD",X"E0",X"7D",X"6A",
		X"C8",X"30",X"27",X"0F",X"AE",X"D4",X"A6",X"11",X"81",X"41",X"27",X"EE",X"81",X"42",X"27",X"EA",
		X"7E",X"11",X"03",X"CC",X"42",X"FF",X"BD",X"E0",X"66",X"86",X"03",X"BD",X"E0",X"7D",X"20",X"F0",
		X"34",X"02",X"A6",X"80",X"1E",X"12",X"BD",X"06",X"43",X"1E",X"12",X"5A",X"26",X"F4",X"35",X"82",
		X"8E",X"CC",X"00",X"6F",X"80",X"8C",X"D0",X"00",X"26",X"F9",X"39",X"34",X"36",X"8E",X"01",X"52",
		X"10",X"8E",X"CC",X"00",X"C6",X"13",X"8D",X"D8",X"35",X"B6",X"34",X"36",X"8E",X"01",X"65",X"10",
		X"8E",X"CC",X"26",X"C6",X"34",X"8D",X"C9",X"BD",X"02",X"50",X"8E",X"CC",X"90",X"BD",X"06",X"43",
		X"35",X"B6",X"50",X"05",X"01",X"03",X"01",X"04",X"01",X"01",X"00",X"00",X"05",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"1A",X"1C",X"0F",X"1D",
		X"0F",X"18",X"1E",X"0F",X"0E",X"0A",X"0C",X"23",X"2D",X"0A",X"0A",X"0A",X"0A",X"0A",X"21",X"13",
		X"16",X"16",X"13",X"0B",X"17",X"1D",X"0A",X"0F",X"16",X"0F",X"0D",X"1E",X"1C",X"19",X"18",X"13",
		X"0D",X"1D",X"0A",X"13",X"18",X"0D",X"2E",X"25",X"29",X"BD",X"02",X"37",X"BD",X"06",X"09",X"B6",
		X"C9",X"80",X"85",X"02",X"26",X"F9",X"B6",X"CC",X"1D",X"84",X"0F",X"27",X"11",X"7F",X"CC",X"1D",
		X"BD",X"02",X"37",X"BD",X"06",X"09",X"BD",X"02",X"DD",X"86",X"40",X"BD",X"F0",X"63",X"B6",X"CC",
		X"1F",X"84",X"0F",X"27",X"0D",X"7F",X"CC",X"1F",X"8D",X"6D",X"BD",X"00",X"12",X"86",X"40",X"BD",
		X"F0",X"63",X"B6",X"CC",X"23",X"84",X"0F",X"27",X"1E",X"7F",X"CC",X"23",X"8D",X"59",X"BD",X"06",
		X"09",X"86",X"09",X"BD",X"E0",X"33",X"BD",X"0A",X"B5",X"86",X"20",X"BD",X"F0",X"63",X"BD",X"02",
		X"50",X"8E",X"CC",X"90",X"BD",X"06",X"43",X"B6",X"CC",X"25",X"84",X"0F",X"27",X"13",X"7F",X"CC",
		X"25",X"8D",X"34",X"BD",X"06",X"09",X"86",X"0F",X"BD",X"E0",X"33",X"BD",X"08",X"E1",X"BD",X"04",
		X"D5",X"B6",X"CC",X"21",X"84",X"0F",X"27",X"0A",X"7F",X"CC",X"21",X"8D",X"1A",X"8D",X"07",X"7E",
		X"F0",X"06",X"8D",X"02",X"20",X"51",X"B6",X"CC",X"1B",X"84",X"0F",X"27",X"09",X"7C",X"CC",X"8E",
		X"7C",X"CC",X"8E",X"7F",X"CC",X"1B",X"39",X"34",X"12",X"8D",X"08",X"8E",X"CC",X"8E",X"BD",X"06",
		X"43",X"35",X"92",X"34",X"34",X"8E",X"CC",X"00",X"10",X"8E",X"CC",X"26",X"8D",X"09",X"35",X"B4",
		X"8E",X"CC",X"26",X"10",X"8E",X"CC",X"8E",X"10",X"9F",X"C5",X"4F",X"E6",X"80",X"C4",X"0F",X"34",
		X"04",X"AB",X"E0",X"9C",X"C5",X"26",X"F4",X"8B",X"37",X"39",X"8D",X"D7",X"34",X"02",X"8E",X"CC",
		X"8E",X"BD",X"06",X"2A",X"A1",X"E0",X"39",X"86",X"90",X"1F",X"8B",X"8D",X"70",X"8D",X"EB",X"27",
		X"3D",X"86",X"14",X"B7",X"C9",X"00",X"BD",X"01",X"2B",X"86",X"14",X"B7",X"C9",X"00",X"8D",X"A7",
		X"86",X"14",X"B7",X"C9",X"00",X"BD",X"06",X"09",X"86",X"14",X"B7",X"C9",X"00",X"8D",X"28",X"BD",
		X"00",X"15",X"BD",X"00",X"0F",X"8D",X"C3",X"27",X"1A",X"86",X"0A",X"BD",X"E0",X"33",X"86",X"14",
		X"B7",X"C9",X"00",X"B6",X"C9",X"80",X"85",X"02",X"27",X"F4",X"6E",X"9F",X"EF",X"FE",X"BD",X"00",
		X"0F",X"20",X"F7",X"86",X"0B",X"20",X"E4",X"8E",X"CD",X"02",X"C6",X"04",X"A6",X"80",X"84",X"0F",
		X"81",X"09",X"23",X"03",X"5A",X"27",X"06",X"8C",X"CD",X"44",X"26",X"F0",X"39",X"86",X"0C",X"BD",
		X"E0",X"33",X"8E",X"CD",X"02",X"6F",X"80",X"8C",X"CD",X"44",X"26",X"F9",X"39",X"8D",X"05",X"27",
		X"FB",X"7E",X"01",X"3A",X"BD",X"02",X"50",X"34",X"02",X"8E",X"CC",X"90",X"BD",X"06",X"2A",X"A1",
		X"E0",X"39",X"86",X"18",X"97",X"D1",X"86",X"08",X"BD",X"F0",X"63",X"B6",X"C9",X"80",X"85",X"08",
		X"27",X"23",X"0A",X"D1",X"26",X"F0",X"10",X"8E",X"CD",X"44",X"8E",X"03",X"8F",X"C6",X"17",X"BD",
		X"00",X"09",X"BD",X"04",X"D5",X"7F",X"C9",X"82",X"B6",X"C9",X"83",X"8A",X"3C",X"B7",X"C9",X"83",
		X"84",X"F7",X"B7",X"C9",X"83",X"39",X"10",X"8E",X"CD",X"7A",X"C6",X"08",X"BD",X"04",X"FC",X"A8",
		X"26",X"84",X"0F",X"27",X"03",X"5A",X"27",X"0E",X"86",X"14",X"B7",X"C9",X"00",X"31",X"2E",X"10",
		X"8C",X"CF",X"AA",X"25",X"E7",X"39",X"86",X"14",X"B7",X"C9",X"00",X"8E",X"03",X"8F",X"10",X"8E",
		X"CD",X"44",X"C6",X"80",X"BD",X"00",X"09",X"8E",X"04",X"0F",X"10",X"8E",X"CE",X"44",X"C6",X"B3",
		X"BD",X"00",X"09",X"BD",X"04",X"D5",X"10",X"8E",X"CD",X"7A",X"BD",X"04",X"F4",X"86",X"14",X"B7",
		X"C9",X"00",X"31",X"2E",X"10",X"8C",X"CF",X"AA",X"25",X"F0",X"86",X"0D",X"7E",X"E0",X"33",X"21",
		X"13",X"16",X"16",X"13",X"0B",X"17",X"1D",X"0A",X"13",X"18",X"10",X"0F",X"1C",X"18",X"19",X"0A",
		X"0A",X"0A",X"0A",X"21",X"13",X"16",X"00",X"10",X"22",X"25",X"16",X"19",X"1F",X"00",X"04",X"84",
		X"93",X"16",X"17",X"1A",X"00",X"04",X"71",X"13",X"16",X"17",X"0B",X"00",X"04",X"61",X"75",X"1A",
		X"0B",X"1C",X"00",X"04",X"52",X"22",X"0F",X"14",X"1D",X"00",X"04",X"42",X"10",X"17",X"16",X"0A",
		X"00",X"04",X"31",X"57",X"1A",X"14",X"0F",X"00",X"04",X"29",X"99",X"15",X"14",X"10",X"00",X"04",
		X"10",X"11",X"11",X"21",X"1D",X"00",X"04",X"05",X"23",X"0B",X"0A",X"16",X"00",X"03",X"99",X"09",
		X"1C",X"0E",X"14",X"00",X"03",X"80",X"01",X"1C",X"17",X"11",X"00",X"03",X"72",X"10",X"23",X"0C",
		X"0A",X"00",X"03",X"61",X"91",X"14",X"11",X"16",X"00",X"03",X"51",X"01",X"17",X"21",X"17",X"00",
		X"03",X"42",X"11",X"0E",X"1C",X"23",X"00",X"03",X"35",X"67",X"11",X"16",X"0C",X"00",X"03",X"28",
		X"90",X"14",X"0A",X"16",X"00",X"03",X"19",X"01",X"16",X"14",X"17",X"00",X"03",X"01",X"57",X"15",
		X"1D",X"12",X"00",X"02",X"92",X"30",X"14",X"19",X"0F",X"00",X"02",X"87",X"77",X"11",X"0B",X"1D",
		X"00",X"02",X"79",X"87",X"17",X"0A",X"1D",X"00",X"02",X"69",X"59",X"1A",X"0A",X"19",X"00",X"02",
		X"58",X"88",X"0C",X"0A",X"21",X"00",X"02",X"46",X"75",X"1A",X"20",X"0B",X"00",X"02",X"33",X"10",
		X"1A",X"10",X"24",X"00",X"02",X"29",X"17",X"1A",X"0B",X"1C",X"00",X"02",X"25",X"52",X"0F",X"14",
		X"1D",X"00",X"02",X"05",X"22",X"17",X"16",X"0A",X"00",X"01",X"71",X"57",X"16",X"19",X"1F",X"00",
		X"01",X"65",X"35",X"0E",X"14",X"21",X"00",X"01",X"55",X"05",X"0C",X"1A",X"0E",X"00",X"01",X"43",
		X"15",X"1C",X"0B",X"17",X"00",X"01",X"31",X"09",X"15",X"20",X"0E",X"00",X"01",X"20",X"10",X"14",
		X"0A",X"17",X"00",X"01",X"17",X"55",X"11",X"21",X"21",X"00",X"01",X"05",X"02",X"20",X"0B",X"22",
		X"00",X"00",X"94",X"05",X"1D",X"0A",X"12",X"00",X"00",X"83",X"11",X"0C",X"0B",X"0E",X"00",X"00",
		X"70",X"01",X"0A",X"0A",X"0A",X"00",X"00",X"40",X"00",X"34",X"34",X"8E",X"04",X"C2",X"C6",X"07",
		X"BD",X"00",X"09",X"35",X"B4",X"34",X"02",X"8D",X"05",X"B7",X"CD",X"72",X"35",X"82",X"34",X"10",
		X"8E",X"CD",X"44",X"4F",X"AB",X"84",X"30",X"01",X"8C",X"CD",X"72",X"27",X"F9",X"8C",X"CD",X"7A",
		X"26",X"F2",X"35",X"90",X"34",X"02",X"8D",X"04",X"A7",X"26",X"35",X"82",X"34",X"24",X"C6",X"0E",
		X"4F",X"C1",X"08",X"27",X"02",X"AB",X"A4",X"31",X"21",X"5A",X"26",X"F5",X"35",X"A4",X"86",X"32",
		X"34",X"02",X"10",X"8E",X"CD",X"7A",X"8D",X"E4",X"A8",X"26",X"84",X"0F",X"27",X"0F",X"BD",X"05",
		X"DE",X"7F",X"CD",X"00",X"7F",X"CD",X"01",X"6A",X"E4",X"27",X"12",X"20",X"E9",X"86",X"03",X"C6",
		X"04",X"8D",X"65",X"25",X"E9",X"31",X"2E",X"10",X"8C",X"CF",X"AA",X"25",X"D9",X"35",X"02",X"8E",
		X"04",X"59",X"10",X"8E",X"CF",X"AA",X"C6",X"2A",X"BD",X"00",X"09",X"8D",X"91",X"B8",X"CD",X"72",
		X"84",X"0F",X"27",X"02",X"8D",X"0F",X"10",X"8E",X"CD",X"44",X"86",X"17",X"C6",X"04",X"8D",X"38",
		X"24",X"02",X"8D",X"01",X"39",X"8E",X"CD",X"44",X"86",X"0A",X"BD",X"06",X"43",X"8C",X"CD",X"6C",
		X"25",X"F8",X"8E",X"CD",X"7A",X"10",X"8E",X"CD",X"44",X"86",X"06",X"BD",X"05",X"FE",X"10",X"8E",
		X"CD",X"6C",X"8D",X"7A",X"8E",X"CD",X"80",X"10",X"8E",X"CD",X"72",X"86",X"08",X"8D",X"6F",X"BD",
		X"04",X"D5",X"10",X"8E",X"CD",X"7A",X"20",X"46",X"34",X"16",X"C6",X"14",X"F7",X"C9",X"00",X"1F",
		X"21",X"BD",X"06",X"3B",X"C1",X"0A",X"25",X"32",X"C1",X"24",X"22",X"2E",X"4A",X"26",X"F2",X"A6",
		X"61",X"BD",X"06",X"3B",X"C4",X"0F",X"C1",X"09",X"22",X"20",X"4A",X"BD",X"06",X"3B",X"34",X"04",
		X"C4",X"0F",X"C1",X"09",X"35",X"04",X"22",X"12",X"C4",X"F0",X"C1",X"99",X"22",X"0C",X"4A",X"26",
		X"EA",X"1C",X"FE",X"86",X"14",X"B7",X"C9",X"00",X"35",X"96",X"1A",X"01",X"20",X"F5",X"34",X"36",
		X"30",X"2E",X"8C",X"CF",X"AA",X"24",X"0F",X"86",X"0E",X"8D",X"13",X"31",X"2E",X"30",X"0E",X"86",
		X"14",X"B7",X"C9",X"00",X"20",X"EC",X"BD",X"04",X"C9",X"BD",X"04",X"F4",X"35",X"B6",X"34",X"36",
		X"E6",X"80",X"E7",X"A0",X"4A",X"26",X"F9",X"35",X"B6",X"34",X"76",X"8E",X"00",X"00",X"1F",X"12",
		X"1F",X"10",X"CE",X"90",X"00",X"86",X"14",X"36",X"34",X"36",X"34",X"36",X"34",X"36",X"34",X"B7",
		X"C9",X"00",X"11",X"83",X"90",X"00",X"25",X"EF",X"35",X"F6",X"A6",X"01",X"84",X"0F",X"34",X"02",
		X"A6",X"81",X"48",X"48",X"48",X"48",X"AB",X"E0",X"39",X"8D",X"EF",X"34",X"02",X"8D",X"EB",X"1F",
		X"89",X"35",X"82",X"34",X"02",X"A7",X"01",X"44",X"44",X"44",X"44",X"A7",X"81",X"35",X"82",X"8D",
		X"F2",X"34",X"02",X"1F",X"98",X"8D",X"EC",X"35",X"82",X"34",X"16",X"86",X"01",X"20",X"02",X"34",
		X"16",X"C4",X"0F",X"58",X"34",X"04",X"58",X"EB",X"E0",X"8E",X"CC",X"FC",X"3A",X"8D",X"CC",X"34",
		X"04",X"8D",X"C8",X"34",X"04",X"8D",X"C4",X"34",X"04",X"AB",X"E4",X"19",X"A7",X"E4",X"A6",X"61",
		X"89",X"00",X"19",X"A7",X"61",X"A6",X"62",X"89",X"00",X"19",X"30",X"1A",X"8D",X"B5",X"35",X"04",
		X"35",X"02",X"8D",X"BB",X"35",X"02",X"35",X"96",X"86",X"0E",X"BD",X"E0",X"33",X"0F",X"C5",X"8E",
		X"0E",X"70",X"CC",X"F1",X"22",X"10",X"8E",X"CD",X"44",X"10",X"9C",X"D9",X"26",X"04",X"C6",X"55",
		X"20",X"07",X"10",X"9C",X"DD",X"26",X"02",X"C6",X"66",X"BD",X"E0",X"17",X"86",X"2B",X"BD",X"E0",
		X"09",X"30",X"89",X"03",X"00",X"86",X"15",X"97",X"CB",X"0A",X"CB",X"27",X"1B",X"1E",X"12",X"BD",
		X"00",X"24",X"81",X"0A",X"2E",X"09",X"0D",X"C5",X"26",X"07",X"10",X"9F",X"C5",X"20",X"02",X"0F",
		X"C5",X"1E",X"12",X"BD",X"E0",X"09",X"20",X"E1",X"0D",X"C5",X"27",X"02",X"9E",X"C5",X"86",X"04",
		X"97",X"CB",X"10",X"8E",X"CD",X"72",X"1E",X"12",X"BD",X"00",X"24",X"1E",X"12",X"8A",X"F0",X"85",
		X"0F",X"26",X"02",X"8A",X"0F",X"BD",X"E0",X"17",X"0A",X"CB",X"1E",X"12",X"BD",X"00",X"24",X"1E",
		X"12",X"BD",X"E0",X"17",X"0A",X"CB",X"26",X"F2",X"8E",X"10",X"80",X"C6",X"33",X"CE",X"E0",X"2C",
		X"DF",X"CE",X"CE",X"E0",X"1E",X"86",X"0D",X"97",X"CB",X"86",X"02",X"97",X"D1",X"86",X"07",X"97",
		X"D0",X"86",X"0F",X"97",X"D6",X"8D",X"48",X"8E",X"3A",X"80",X"86",X"0D",X"97",X"CB",X"86",X"15",
		X"97",X"D1",X"8D",X"3B",X"8E",X"64",X"80",X"86",X"0D",X"97",X"CB",X"86",X"28",X"97",X"D1",X"8D",
		X"2E",X"8E",X"13",X"36",X"10",X"8E",X"CF",X"AA",X"C6",X"11",X"CE",X"E0",X"17",X"DF",X"CE",X"CE",
		X"E0",X"09",X"86",X"03",X"97",X"CB",X"86",X"01",X"97",X"D1",X"86",X"0A",X"97",X"D0",X"86",X"15",
		X"97",X"D6",X"8D",X"0B",X"8E",X"53",X"36",X"86",X"03",X"97",X"CB",X"86",X"04",X"97",X"D1",X"9F",
		X"C8",X"34",X"04",X"C6",X"03",X"D7",X"D8",X"5C",X"D7",X"D5",X"E6",X"E4",X"10",X"9C",X"D9",X"27",
		X"05",X"10",X"9C",X"DB",X"26",X"02",X"C6",X"55",X"10",X"9C",X"DD",X"27",X"05",X"10",X"9C",X"DF",
		X"26",X"02",X"C6",X"66",X"96",X"D1",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"AD",X"9F",X"90",X"CE",
		X"86",X"2B",X"AD",X"C4",X"86",X"0A",X"AD",X"C4",X"1E",X"12",X"BD",X"00",X"24",X"1E",X"12",X"AD",
		X"C4",X"0A",X"D8",X"26",X"F3",X"9F",X"C5",X"9E",X"C8",X"1E",X"01",X"D6",X"C6",X"9B",X"D6",X"1E",
		X"01",X"0F",X"CC",X"1E",X"12",X"BD",X"00",X"24",X"1E",X"12",X"0D",X"CC",X"26",X"1A",X"34",X"02",
		X"86",X"04",X"91",X"D5",X"26",X"04",X"35",X"02",X"20",X"06",X"35",X"02",X"85",X"F0",X"26",X"08",
		X"8A",X"F0",X"85",X"0F",X"26",X"02",X"8A",X"0F",X"97",X"CC",X"03",X"CC",X"AD",X"9F",X"90",X"CE",
		X"0A",X"D5",X"26",X"CF",X"9F",X"C5",X"9E",X"C8",X"1E",X"01",X"D6",X"C6",X"DB",X"D0",X"1E",X"01",
		X"96",X"D1",X"8B",X"01",X"19",X"97",X"D1",X"0A",X"CB",X"35",X"04",X"10",X"26",X"FF",X"62",X"39",
		X"34",X"12",X"9B",X"E1",X"19",X"24",X"02",X"86",X"99",X"97",X"E1",X"8E",X"CD",X"00",X"BD",X"06",
		X"43",X"35",X"12",X"7E",X"11",X"06",X"34",X"16",X"C6",X"03",X"20",X"0A",X"34",X"16",X"C6",X"02",
		X"20",X"04",X"34",X"16",X"C6",X"01",X"BD",X"06",X"59",X"58",X"8E",X"CC",X"06",X"3A",X"BD",X"06",
		X"3B",X"8D",X"62",X"96",X"E3",X"34",X"04",X"AB",X"E4",X"97",X"E3",X"96",X"E2",X"AB",X"E0",X"97",
		X"E2",X"8E",X"CC",X"12",X"BD",X"06",X"3B",X"8D",X"4C",X"34",X"04",X"A1",X"E0",X"24",X"02",X"35",
		X"96",X"8E",X"CC",X"0E",X"BD",X"06",X"3B",X"8D",X"3C",X"8D",X"24",X"34",X"02",X"D7",X"E2",X"8E",
		X"CC",X"10",X"BD",X"06",X"3B",X"96",X"E3",X"8D",X"2C",X"8D",X"14",X"4D",X"27",X"04",X"0F",X"E2",
		X"0F",X"E3",X"AB",X"E0",X"19",X"C6",X"04",X"BD",X"06",X"5F",X"BD",X"08",X"20",X"35",X"96",X"34",
		X"04",X"5D",X"26",X"03",X"4F",X"35",X"84",X"1E",X"89",X"86",X"99",X"8B",X"01",X"19",X"E0",X"E4",
		X"24",X"F9",X"EB",X"E0",X"39",X"34",X"02",X"4F",X"C1",X"10",X"25",X"06",X"8B",X"0A",X"C0",X"10",
		X"20",X"F6",X"34",X"04",X"AB",X"E0",X"1F",X"89",X"35",X"82",X"34",X"04",X"1F",X"89",X"4F",X"C1",
		X"0A",X"25",X"07",X"8B",X"10",X"19",X"C0",X"0A",X"20",X"F5",X"34",X"04",X"AB",X"E0",X"19",X"35",
		X"84",X"CE",X"B0",X"00",X"8E",X"CC",X"16",X"BD",X"06",X"3B",X"8D",X"C9",X"E7",X"42",X"CC",X"0A",
		X"25",X"BD",X"09",X"1B",X"8E",X"20",X"80",X"AF",X"49",X"CC",X"00",X"63",X"ED",X"46",X"86",X"77",
		X"A7",X"48",X"BD",X"0A",X"29",X"BD",X"09",X"38",X"24",X"F8",X"C6",X"14",X"8E",X"CD",X"44",X"31",
		X"C8",X"11",X"A6",X"A0",X"BD",X"06",X"43",X"5A",X"26",X"F8",X"39",X"34",X"16",X"A7",X"44",X"E7",
		X"45",X"86",X"0A",X"A7",X"C8",X"10",X"A7",X"4F",X"6F",X"43",X"30",X"C8",X"11",X"C6",X"19",X"86",
		X"0A",X"A7",X"80",X"5A",X"26",X"FB",X"35",X"96",X"4F",X"E6",X"43",X"27",X"0E",X"34",X"04",X"CB",
		X"10",X"E6",X"C5",X"BD",X"E0",X"5D",X"35",X"04",X"5A",X"26",X"F2",X"AE",X"49",X"30",X"8B",X"AF",
		X"4B",X"C6",X"11",X"EB",X"43",X"A6",X"C5",X"BD",X"09",X"E1",X"AD",X"D8",X"06",X"C4",X"FF",X"26",
		X"09",X"6F",X"4F",X"C6",X"0A",X"E7",X"C8",X"10",X"20",X"5D",X"6D",X"4F",X"27",X"04",X"6A",X"4F",
		X"20",X"55",X"34",X"06",X"A6",X"C8",X"10",X"81",X"04",X"23",X"02",X"80",X"02",X"A7",X"C8",X"10",
		X"A7",X"4F",X"35",X"06",X"C5",X"30",X"27",X"0F",X"81",X"25",X"27",X"2D",X"8D",X"4E",X"6C",X"43",
		X"6A",X"42",X"26",X"33",X"1A",X"01",X"39",X"C5",X"03",X"27",X"0D",X"8D",X"3C",X"A1",X"45",X"26",
		X"04",X"A6",X"44",X"20",X"22",X"4C",X"20",X"1F",X"C5",X"0C",X"27",X"0D",X"8D",X"2B",X"A1",X"44",
		X"26",X"04",X"A6",X"45",X"20",X"11",X"4A",X"20",X"0E",X"6D",X"43",X"27",X"0A",X"8D",X"1A",X"8D",
		X"1B",X"6C",X"42",X"6A",X"43",X"20",X"02",X"8D",X"03",X"1C",X"FE",X"39",X"C6",X"11",X"EB",X"43",
		X"A7",X"C5",X"E6",X"48",X"AE",X"4B",X"7E",X"E0",X"09",X"5F",X"20",X"F8",X"34",X"27",X"5F",X"20",
		X"04",X"34",X"27",X"E6",X"48",X"1A",X"F0",X"F7",X"C8",X"81",X"CC",X"0A",X"21",X"FD",X"C8",X"82",
		X"AE",X"4B",X"30",X"08",X"CC",X"04",X"02",X"8D",X"19",X"CC",X"0A",X"22",X"FD",X"C8",X"82",X"E6",
		X"42",X"5A",X"2F",X"0C",X"4F",X"1F",X"02",X"CC",X"03",X"01",X"8D",X"06",X"31",X"3F",X"26",X"F7",
		X"35",X"A7",X"FD",X"C8",X"86",X"BF",X"C8",X"84",X"C6",X"1A",X"F7",X"C8",X"80",X"5F",X"30",X"8B",
		X"39",X"11",X"11",X"11",X"10",X"11",X"11",X"11",X"10",X"34",X"16",X"86",X"04",X"BD",X"F0",X"63",
		X"35",X"96",X"C6",X"66",X"D7",X"D8",X"C6",X"CA",X"8D",X"04",X"C6",X"D8",X"20",X"2C",X"34",X"76",
		X"8E",X"CC",X"8A",X"BD",X"00",X"24",X"1F",X"02",X"1F",X"03",X"8E",X"CC",X"26",X"D6",X"D8",X"BD",
		X"00",X"24",X"1E",X"12",X"81",X"0A",X"27",X"02",X"1F",X"13",X"BD",X"E0",X"09",X"1E",X"12",X"8C",
		X"CC",X"58",X"26",X"EB",X"11",X"83",X"8E",X"00",X"35",X"F6",X"34",X"76",X"8E",X"CC",X"8C",X"BD",
		X"00",X"24",X"1F",X"02",X"8E",X"CC",X"58",X"D6",X"D8",X"BD",X"00",X"24",X"1E",X"12",X"81",X"0A",
		X"27",X"02",X"1F",X"13",X"BD",X"E0",X"09",X"1E",X"12",X"8C",X"CC",X"8A",X"26",X"EB",X"11",X"83",
		X"8E",X"00",X"35",X"F6",X"CE",X"B0",X"00",X"AF",X"49",X"CC",X"00",X"34",X"BD",X"09",X"1B",X"C6",
		X"19",X"E7",X"42",X"CC",X"00",X"63",X"ED",X"46",X"86",X"77",X"A7",X"48",X"BD",X"0A",X"29",X"BD",
		X"09",X"38",X"24",X"F8",X"39",X"8E",X"25",X"60",X"8D",X"DA",X"C6",X"19",X"8E",X"CC",X"26",X"31",
		X"C8",X"11",X"A6",X"A0",X"BD",X"06",X"43",X"5A",X"26",X"F8",X"86",X"25",X"8E",X"CC",X"8A",X"BD",
		X"06",X"43",X"C6",X"88",X"8D",X"2F",X"86",X"34",X"C6",X"22",X"8E",X"48",X"6A",X"BD",X"E0",X"09",
		X"CE",X"0B",X"15",X"8E",X"CC",X"8A",X"BD",X"0B",X"72",X"C6",X"60",X"BD",X"0A",X"3E",X"25",X"04",
		X"91",X"E8",X"25",X"08",X"96",X"E8",X"8E",X"CC",X"8A",X"BD",X"06",X"43",X"86",X"22",X"97",X"D8",
		X"BD",X"0A",X"3E",X"20",X"DE",X"86",X"4E",X"8E",X"25",X"90",X"BD",X"E0",X"10",X"86",X"4F",X"8E",
		X"25",X"A0",X"7E",X"E0",X"10",X"86",X"34",X"C6",X"00",X"8E",X"48",X"6A",X"BD",X"E0",X"09",X"8D",
		X"E4",X"8E",X"25",X"70",X"BD",X"0A",X"94",X"C6",X"19",X"8E",X"CC",X"58",X"31",X"C8",X"11",X"A6",
		X"A0",X"BD",X"06",X"43",X"5A",X"26",X"F8",X"86",X"25",X"8E",X"CC",X"8C",X"BD",X"06",X"43",X"C6",
		X"88",X"8D",X"C2",X"86",X"34",X"C6",X"22",X"8E",X"48",X"7A",X"BD",X"E0",X"09",X"CE",X"0B",X"71",
		X"8E",X"CC",X"8C",X"8D",X"1D",X"C6",X"70",X"BD",X"0A",X"6A",X"25",X"04",X"91",X"E8",X"25",X"08",
		X"96",X"E8",X"8E",X"CC",X"8C",X"BD",X"06",X"43",X"86",X"22",X"97",X"D8",X"BD",X"0A",X"6A",X"20",
		X"DF",X"39",X"F6",X"C9",X"80",X"C5",X"02",X"27",X"04",X"32",X"62",X"6E",X"C4",X"BD",X"0A",X"29",
		X"BD",X"00",X"63",X"C4",X"F0",X"27",X"EB",X"0F",X"F2",X"0F",X"F3",X"BD",X"06",X"2A",X"97",X"C0",
		X"C5",X"5F",X"26",X"07",X"81",X"08",X"23",X"DA",X"4A",X"20",X"01",X"4C",X"97",X"E8",X"0F",X"D8",
		X"96",X"C0",X"39",X"A6",X"84",X"84",X"F0",X"27",X"07",X"CC",X"99",X"99",X"ED",X"81",X"ED",X"81",
		X"39",X"0F",X"E4",X"4F",X"5F",X"DD",X"D9",X"DD",X"DB",X"DD",X"DD",X"DD",X"DF",X"B6",X"CC",X"05",
		X"44",X"25",X"03",X"7E",X"11",X"03",X"8E",X"90",X"2B",X"8D",X"D8",X"8E",X"90",X"3A",X"8D",X"D3",
		X"0D",X"49",X"27",X"5B",X"8E",X"90",X"2B",X"10",X"8E",X"90",X"3A",X"BD",X"0F",X"04",X"25",X"4F",
		X"1E",X"21",X"BD",X"0E",X"C8",X"24",X"23",X"0C",X"E4",X"10",X"8E",X"0E",X"51",X"86",X"42",X"5F",
		X"BD",X"E0",X"63",X"86",X"10",X"A7",X"33",X"86",X"01",X"A7",X"A8",X"2F",X"8E",X"90",X"3A",X"AF",
		X"A8",X"2B",X"8E",X"70",X"A0",X"AF",X"A8",X"2D",X"20",X"12",X"8E",X"90",X"3A",X"AF",X"C8",X"2B",
		X"8E",X"70",X"A0",X"AF",X"C8",X"2D",X"86",X"01",X"C6",X"42",X"8D",X"67",X"8E",X"90",X"2B",X"AF",
		X"C8",X"2B",X"8E",X"20",X"A0",X"AF",X"C8",X"2D",X"4F",X"C6",X"41",X"8D",X"56",X"20",X"51",X"8E",
		X"90",X"2B",X"BD",X"0E",X"C8",X"24",X"22",X"0C",X"E4",X"10",X"8E",X"0E",X"51",X"86",X"42",X"5F",
		X"BD",X"E0",X"63",X"86",X"10",X"A7",X"33",X"4F",X"A7",X"A8",X"2F",X"8E",X"90",X"2B",X"AF",X"A8",
		X"2B",X"8E",X"20",X"A0",X"AF",X"A8",X"2D",X"20",X"11",X"8E",X"90",X"2B",X"AF",X"C8",X"2B",X"8E",
		X"20",X"A0",X"AF",X"C8",X"2D",X"4F",X"C6",X"42",X"8D",X"19",X"0D",X"49",X"27",X"12",X"8E",X"90",
		X"3A",X"AF",X"C8",X"2B",X"8E",X"70",X"A0",X"AF",X"C8",X"2D",X"86",X"01",X"C6",X"41",X"8D",X"03",
		X"7E",X"00",X"BE",X"BD",X"0E",X"CE",X"24",X"24",X"0C",X"E4",X"34",X"02",X"10",X"8E",X"0C",X"D5",
		X"1F",X"98",X"5F",X"BD",X"E0",X"63",X"86",X"10",X"A7",X"33",X"35",X"02",X"A7",X"A8",X"2F",X"AE",
		X"C8",X"2B",X"AF",X"A8",X"2B",X"AE",X"C8",X"2D",X"AF",X"A8",X"2D",X"39",X"BD",X"0E",X"EB",X"24",
		X"23",X"0C",X"E4",X"34",X"02",X"10",X"8E",X"0C",X"D5",X"1F",X"98",X"5F",X"BD",X"E0",X"63",X"86",
		X"08",X"A7",X"33",X"35",X"02",X"A7",X"A8",X"2F",X"AE",X"C8",X"2B",X"AF",X"A8",X"2B",X"AE",X"C8",
		X"2D",X"AF",X"A8",X"2D",X"39",X"6F",X"C8",X"2A",X"E6",X"C8",X"2F",X"26",X"0E",X"8E",X"0A",X"B0",
		X"CC",X"00",X"63",X"ED",X"46",X"34",X"04",X"C6",X"55",X"20",X"0A",X"8E",X"58",X"B0",X"CC",X"00",
		X"6F",X"ED",X"46",X"C6",X"66",X"86",X"54",X"BD",X"E0",X"10",X"1F",X"98",X"8E",X"0D",X"07",X"AF",
		X"4D",X"AE",X"C8",X"2D",X"7E",X"0F",X"3C",X"A6",X"51",X"81",X"42",X"27",X"1F",X"ED",X"C8",X"30",
		X"AF",X"C8",X"32",X"10",X"AF",X"42",X"86",X"01",X"BD",X"E0",X"7D",X"AE",X"C4",X"A6",X"11",X"81",
		X"42",X"27",X"F3",X"EC",X"C8",X"30",X"AE",X"C8",X"32",X"10",X"AE",X"42",X"BD",X"0E",X"CE",X"24",
		X"13",X"6D",X"C8",X"2F",X"26",X"05",X"10",X"9F",X"DB",X"20",X"03",X"10",X"9F",X"DF",X"8E",X"CF",
		X"F0",X"BD",X"0E",X"1F",X"BD",X"0E",X"EB",X"24",X"18",X"6D",X"C8",X"2A",X"27",X"1C",X"30",X"C8",
		X"11",X"10",X"8E",X"CD",X"6C",X"C6",X"03",X"BD",X"01",X"10",X"BD",X"04",X"D5",X"86",X"05",X"8D",
		X"74",X"24",X"6F",X"1F",X"12",X"BD",X"05",X"DE",X"20",X"50",X"30",X"A9",X"32",X"9A",X"26",X"2B",
		X"8E",X"CF",X"9C",X"BD",X"0E",X"3B",X"31",X"26",X"AE",X"C8",X"2B",X"C6",X"04",X"BD",X"01",X"10",
		X"10",X"8E",X"CD",X"44",X"6D",X"C8",X"2F",X"26",X"05",X"10",X"9F",X"D9",X"20",X"03",X"10",X"9F",
		X"DD",X"30",X"C8",X"11",X"C6",X"14",X"BD",X"01",X"10",X"20",X"B3",X"BD",X"0D",X"D9",X"34",X"01",
		X"34",X"10",X"10",X"AC",X"E1",X"22",X"0F",X"8D",X"76",X"6D",X"C8",X"2F",X"26",X"05",X"10",X"9F",
		X"D9",X"20",X"03",X"10",X"9F",X"DD",X"35",X"01",X"24",X"18",X"8E",X"90",X"D9",X"31",X"C4",X"AE",
		X"C8",X"2D",X"30",X"89",X"EA",X"F6",X"86",X"56",X"E6",X"48",X"BD",X"E0",X"10",X"86",X"60",X"BD",
		X"E0",X"7D",X"7E",X"E0",X"69",X"34",X"26",X"20",X"0C",X"34",X"26",X"8E",X"CD",X"6C",X"8D",X"24",
		X"86",X"04",X"25",X"01",X"4C",X"97",X"C5",X"8E",X"CD",X"7A",X"8D",X"18",X"24",X"04",X"0A",X"C5",
		X"27",X"0E",X"30",X"0E",X"8C",X"CF",X"AA",X"25",X"F1",X"8E",X"CF",X"9C",X"1C",X"FE",X"35",X"A6",
		X"1A",X"01",X"35",X"A6",X"34",X"10",X"31",X"C4",X"31",X"C8",X"11",X"C6",X"03",X"BD",X"06",X"2A",
		X"A1",X"A0",X"26",X"07",X"5A",X"26",X"F6",X"1A",X"01",X"35",X"90",X"1C",X"FE",X"35",X"90",X"34",
		X"20",X"BD",X"0E",X"3B",X"30",X"C4",X"30",X"C8",X"11",X"C6",X"03",X"BD",X"01",X"10",X"AE",X"C8",
		X"2B",X"C6",X"04",X"BD",X"01",X"10",X"35",X"20",X"7E",X"04",X"F4",X"34",X"30",X"1F",X"12",X"10",
		X"AC",X"62",X"27",X"0B",X"30",X"32",X"86",X"0E",X"BD",X"05",X"FE",X"31",X"32",X"20",X"F0",X"35",
		X"B0",X"86",X"FF",X"A7",X"C8",X"2A",X"31",X"C4",X"A6",X"C8",X"2F",X"26",X"09",X"CC",X"00",X"63",
		X"ED",X"46",X"C6",X"55",X"20",X"07",X"CC",X"00",X"6F",X"ED",X"46",X"C6",X"66",X"86",X"53",X"8E",
		X"1E",X"5B",X"BD",X"E0",X"10",X"1F",X"98",X"8E",X"0E",X"7F",X"AF",X"4D",X"7E",X"0F",X"2E",X"30",
		X"C8",X"11",X"10",X"8E",X"CD",X"44",X"C6",X"14",X"BD",X"01",X"10",X"10",X"8E",X"CD",X"6C",X"8E",
		X"CF",X"9C",X"BD",X"0E",X"3B",X"10",X"8E",X"CD",X"7A",X"BD",X"04",X"F4",X"AE",X"C8",X"2B",X"10",
		X"8E",X"CD",X"72",X"C6",X"04",X"BD",X"01",X"10",X"8E",X"04",X"C2",X"10",X"8E",X"CD",X"6C",X"C6",
		X"03",X"BD",X"01",X"10",X"BD",X"04",X"D5",X"8E",X"CD",X"44",X"A6",X"C8",X"2F",X"26",X"04",X"9F",
		X"D9",X"20",X"02",X"9F",X"DD",X"7E",X"0C",X"D8",X"10",X"8E",X"CD",X"72",X"20",X"36",X"34",X"16",
		X"10",X"8E",X"CF",X"B0",X"AE",X"C8",X"2B",X"8D",X"2B",X"25",X"0C",X"31",X"2E",X"10",X"8C",X"CF",
		X"FE",X"25",X"F4",X"1C",X"FE",X"35",X"96",X"31",X"3A",X"35",X"96",X"34",X"16",X"10",X"8E",X"CD",
		X"72",X"AE",X"C8",X"2B",X"8D",X"0E",X"25",X"EF",X"31",X"2E",X"10",X"8C",X"CF",X"9C",X"25",X"F4",
		X"1C",X"FE",X"35",X"96",X"34",X"36",X"1E",X"12",X"C6",X"04",X"8D",X"17",X"C1",X"04",X"26",X"02",
		X"84",X"0F",X"A1",X"A0",X"22",X"05",X"25",X"07",X"5A",X"26",X"EF",X"1C",X"FE",X"35",X"B6",X"1A",
		X"01",X"35",X"B6",X"8C",X"C0",X"00",X"25",X"03",X"7E",X"06",X"2A",X"A6",X"80",X"39",X"8E",X"CC",
		X"16",X"BD",X"06",X"3B",X"BD",X"08",X"B5",X"8E",X"26",X"43",X"20",X"02",X"C6",X"03",X"A7",X"48",
		X"E7",X"42",X"AF",X"49",X"CC",X"0A",X"25",X"BD",X"09",X"1B",X"86",X"01",X"BD",X"E0",X"7D",X"BD",
		X"09",X"38",X"24",X"F6",X"6E",X"D8",X"0D",X"FC",X"0F",X"D4",X"8D",X"53",X"8D",X"2A",X"8E",X"0F",
		X"D4",X"EC",X"81",X"9F",X"C5",X"8D",X"48",X"86",X"80",X"97",X"E8",X"4F",X"BD",X"F0",X"63",X"BD",
		X"F0",X"6C",X"25",X"13",X"B6",X"C9",X"80",X"46",X"24",X"F1",X"0A",X"E8",X"26",X"ED",X"9E",X"C5",
		X"8C",X"0F",X"FC",X"25",X"DC",X"20",X"D7",X"39",X"8E",X"00",X"00",X"10",X"8E",X"0F",X"FC",X"9F",
		X"C5",X"30",X"89",X"09",X"00",X"A6",X"A0",X"1F",X"89",X"ED",X"83",X"C6",X"14",X"F7",X"C9",X"00",
		X"9C",X"C5",X"26",X"F3",X"30",X"89",X"09",X"00",X"10",X"8C",X"10",X"0C",X"26",X"E1",X"39",X"34",
		X"06",X"8E",X"86",X"20",X"B6",X"BF",X"FF",X"34",X"02",X"86",X"03",X"B7",X"BF",X"FF",X"B7",X"C8",
		X"00",X"EC",X"61",X"ED",X"81",X"8C",X"86",X"40",X"25",X"F9",X"35",X"02",X"B7",X"BF",X"FF",X"B7",
		X"C8",X"00",X"35",X"86",X"00",X"F1",X"00",X"F2",X"00",X"F4",X"00",X"F8",X"00",X"FF",X"01",X"F0",
		X"02",X"F0",X"04",X"F0",X"08",X"F0",X"0F",X"F0",X"10",X"F0",X"20",X"F0",X"40",X"F0",X"80",X"F0",
		X"F0",X"F0",X"FF",X"1F",X"FF",X"2F",X"FF",X"4F",X"FF",X"8F",X"FF",X"FF",X"FF",X"11",X"EE",X"22",
		X"DD",X"33",X"CC",X"44",X"BB",X"55",X"AA",X"66",X"99",X"77",X"88",X"FF",X"20",X"49",X"4E",X"46",
		X"45",X"52",X"4E",X"4F",X"20",X"2D",X"20",X"28",X"43",X"29",X"31",X"39",X"38",X"34",X"20",X"57",
		X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",
		X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"1C",X"1E",X"7E",X"1C",X"44",X"7E",X"25",X"51",X"29",X"85",X"7E",X"1C",X"70",X"7E",X"25",
		X"59",X"24",X"64",X"12",X"8C",X"12",X"CA",X"7E",X"13",X"08",X"7E",X"16",X"84",X"7E",X"11",X"E6",
		X"7E",X"11",X"9E",X"7E",X"16",X"33",X"7E",X"13",X"E9",X"7E",X"14",X"0A",X"7E",X"1C",X"22",X"7E",
		X"11",X"CF",X"7E",X"1C",X"05",X"7E",X"11",X"4B",X"7E",X"1E",X"4D",X"7E",X"25",X"8C",X"7E",X"27",
		X"47",X"7E",X"25",X"6F",X"7E",X"16",X"7F",X"18",X"EA",X"19",X"33",X"6F",X"E2",X"6F",X"E2",X"6F",
		X"E2",X"6F",X"E2",X"C5",X"0F",X"27",X"06",X"8D",X"27",X"C5",X"0F",X"27",X"FA",X"C5",X"F0",X"27",
		X"14",X"86",X"04",X"54",X"68",X"23",X"69",X"22",X"69",X"21",X"69",X"A4",X"4A",X"26",X"F4",X"8D",
		X"0F",X"C5",X"0F",X"26",X"FA",X"6F",X"A4",X"35",X"06",X"ED",X"21",X"35",X"06",X"A7",X"23",X"39",
		X"A6",X"23",X"AB",X"65",X"19",X"A7",X"65",X"A6",X"22",X"A9",X"64",X"19",X"A7",X"64",X"A6",X"21",
		X"A9",X"63",X"19",X"A7",X"63",X"A6",X"A4",X"A9",X"62",X"19",X"A7",X"62",X"5A",X"39",X"8E",X"90",
		X"90",X"4F",X"5F",X"A7",X"80",X"8C",X"90",X"B6",X"25",X"F9",X"8E",X"B7",X"16",X"A7",X"80",X"8C",
		X"B8",X"3B",X"25",X"F9",X"DD",X"36",X"DD",X"38",X"DD",X"45",X"DD",X"47",X"0C",X"2F",X"0C",X"3E",
		X"BD",X"E0",X"AA",X"BD",X"11",X"CF",X"BD",X"00",X"21",X"BE",X"E0",X"7B",X"7E",X"E0",X"6F",X"34",
		X"16",X"CC",X"00",X"00",X"8E",X"C0",X"00",X"ED",X"81",X"ED",X"81",X"ED",X"81",X"ED",X"81",X"8C",
		X"C8",X"00",X"25",X"F3",X"35",X"96",X"34",X"76",X"0F",X"BB",X"0F",X"BC",X"0F",X"BD",X"0F",X"BE",
		X"AE",X"C8",X"22",X"10",X"AE",X"88",X"14",X"2A",X"1D",X"50",X"CB",X"07",X"8E",X"90",X"BB",X"54",
		X"3A",X"25",X"0C",X"1F",X"89",X"48",X"48",X"48",X"48",X"54",X"54",X"54",X"54",X"E7",X"1F",X"A7",
		X"84",X"AE",X"C8",X"22",X"8D",X"02",X"35",X"F6",X"96",X"BE",X"AB",X"23",X"19",X"A7",X"23",X"96",
		X"BD",X"A9",X"22",X"19",X"A7",X"22",X"96",X"BC",X"A9",X"21",X"19",X"A7",X"21",X"96",X"BB",X"A9",
		X"A4",X"19",X"24",X"02",X"8B",X"10",X"A7",X"A4",X"96",X"BE",X"AB",X"2E",X"19",X"A7",X"2E",X"96",
		X"BD",X"A9",X"2D",X"19",X"A7",X"2D",X"96",X"BC",X"A9",X"2C",X"19",X"A7",X"2C",X"96",X"BB",X"A9",
		X"2B",X"19",X"24",X"02",X"8B",X"10",X"A7",X"2B",X"6C",X"24",X"DC",X"69",X"27",X"2D",X"EC",X"21",
		X"AB",X"28",X"19",X"10",X"A3",X"29",X"25",X"23",X"A6",X"2A",X"9B",X"6A",X"19",X"A7",X"2A",X"A6",
		X"29",X"99",X"69",X"19",X"A7",X"29",X"81",X"30",X"25",X"0C",X"8B",X"80",X"19",X"A7",X"29",X"A6",
		X"28",X"8B",X"80",X"19",X"A7",X"28",X"BD",X"13",X"E9",X"20",X"D3",X"39",X"90",X"2F",X"1A",X"55",
		X"90",X"2B",X"0A",X"11",X"13",X"6E",X"90",X"2C",X"0D",X"11",X"13",X"6A",X"90",X"2C",X"10",X"11",
		X"13",X"6E",X"90",X"2D",X"13",X"11",X"13",X"6A",X"90",X"2D",X"16",X"11",X"13",X"6E",X"90",X"2E",
		X"19",X"11",X"13",X"6A",X"90",X"2E",X"1C",X"11",X"13",X"6E",X"90",X"30",X"0E",X"1A",X"13",X"79",
		X"90",X"32",X"1D",X"1A",X"13",X"7E",X"00",X"00",X"00",X"00",X"90",X"3E",X"1A",X"66",X"90",X"3A",
		X"71",X"11",X"13",X"6E",X"90",X"3B",X"74",X"11",X"13",X"6A",X"90",X"3B",X"77",X"11",X"13",X"6E",
		X"90",X"3C",X"7A",X"11",X"13",X"6A",X"90",X"3C",X"7D",X"11",X"13",X"6E",X"90",X"3D",X"80",X"11",
		X"13",X"6A",X"90",X"3D",X"83",X"11",X"13",X"6E",X"90",X"3F",X"75",X"1A",X"13",X"74",X"90",X"41",
		X"84",X"1A",X"13",X"7E",X"00",X"00",X"00",X"00",X"AE",X"48",X"20",X"2E",X"AF",X"4A",X"10",X"AE",
		X"48",X"EE",X"22",X"10",X"AE",X"02",X"27",X"0D",X"E6",X"94",X"AD",X"98",X"04",X"DE",X"21",X"AE",
		X"4A",X"30",X"06",X"20",X"E7",X"DE",X"21",X"86",X"03",X"A7",X"4D",X"86",X"02",X"BD",X"E0",X"7D",
		X"AE",X"48",X"E6",X"94",X"26",X"04",X"6A",X"4D",X"26",X"F1",X"6F",X"94",X"30",X"04",X"E6",X"94",
		X"26",X"CA",X"30",X"06",X"E6",X"94",X"27",X"08",X"C4",X"F0",X"26",X"C0",X"30",X"06",X"20",X"BC",
		X"30",X"0C",X"E6",X"94",X"27",X"08",X"C4",X"F0",X"26",X"B2",X"30",X"06",X"20",X"AE",X"30",X"0C",
		X"E6",X"94",X"C4",X"F0",X"26",X"A6",X"30",X"06",X"20",X"A2",X"56",X"56",X"56",X"56",X"8E",X"30",
		X"00",X"7E",X"E0",X"60",X"8E",X"29",X"76",X"20",X"0B",X"8E",X"29",X"6A",X"20",X"06",X"8E",X"29",
		X"5E",X"CE",X"1A",X"88",X"C1",X"03",X"22",X"2A",X"1A",X"F0",X"EE",X"81",X"FF",X"C8",X"86",X"BF",
		X"C8",X"82",X"7F",X"C8",X"81",X"86",X"02",X"8D",X"07",X"8D",X"05",X"8D",X"03",X"1C",X"EF",X"39",
		X"5D",X"2E",X"02",X"86",X"12",X"5A",X"10",X"BF",X"C8",X"84",X"31",X"A9",X"02",X"00",X"B7",X"C8",
		X"80",X"39",X"34",X"04",X"C5",X"F0",X"26",X"04",X"8D",X"0A",X"20",X"02",X"8D",X"21",X"35",X"04",
		X"8D",X"21",X"20",X"00",X"1A",X"F0",X"8E",X"03",X"05",X"BF",X"C8",X"86",X"10",X"BF",X"C8",X"84",
		X"31",X"A9",X"02",X"00",X"7F",X"C8",X"81",X"86",X"12",X"B7",X"C8",X"80",X"1C",X"EF",X"39",X"56",
		X"56",X"56",X"56",X"8E",X"30",X"6A",X"7E",X"E0",X"60",X"34",X"30",X"8E",X"29",X"82",X"BD",X"E0",
		X"75",X"AE",X"E4",X"AE",X"88",X"14",X"27",X"10",X"A6",X"05",X"8B",X"01",X"19",X"27",X"09",X"A7",
		X"05",X"6C",X"06",X"C6",X"05",X"BD",X"00",X"1E",X"35",X"B0",X"34",X"10",X"AE",X"88",X"14",X"27",
		X"1A",X"A6",X"06",X"27",X"02",X"6A",X"06",X"A6",X"05",X"27",X"10",X"D6",X"68",X"2A",X"05",X"C6",
		X"07",X"BD",X"00",X"1E",X"8B",X"99",X"19",X"A7",X"05",X"86",X"01",X"35",X"90",X"00",X"20",X"00",
		X"20",X"00",X"20",X"00",X"40",X"F6",X"42",X"42",X"14",X"21",X"02",X"00",X"12",X"00",X"0C",X"00",
		X"08",X"00",X"00",X"F6",X"42",X"42",X"14",X"21",X"FE",X"00",X"06",X"00",X"04",X"00",X"02",X"00",
		X"00",X"F6",X"42",X"42",X"14",X"21",X"FE",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"00",X"F6",
		X"42",X"42",X"14",X"21",X"FD",X"00",X"78",X"00",X"50",X"00",X"32",X"00",X"01",X"F2",X"22",X"22",
		X"12",X"21",X"FC",X"00",X"50",X"00",X"3C",X"00",X"28",X"00",X"01",X"F2",X"22",X"22",X"12",X"21",
		X"F8",X"00",X"1E",X"00",X"1E",X"00",X"1E",X"00",X"01",X"F2",X"22",X"22",X"12",X"21",X"F0",X"00",
		X"12",X"00",X"0E",X"00",X"0A",X"00",X"05",X"F6",X"42",X"42",X"14",X"21",X"FC",X"00",X"08",X"00",
		X"06",X"00",X"04",X"00",X"01",X"F6",X"42",X"42",X"14",X"21",X"FC",X"00",X"20",X"00",X"18",X"00",
		X"0C",X"00",X"01",X"F6",X"42",X"42",X"14",X"21",X"FC",X"00",X"30",X"00",X"28",X"00",X"1E",X"00",
		X"01",X"F6",X"42",X"42",X"14",X"21",X"FC",X"00",X"28",X"00",X"20",X"00",X"18",X"00",X"01",X"F6",
		X"42",X"42",X"14",X"21",X"FA",X"00",X"1E",X"00",X"18",X"00",X"12",X"00",X"01",X"F6",X"42",X"42",
		X"14",X"21",X"F8",X"00",X"1E",X"00",X"1E",X"00",X"0F",X"00",X"01",X"F6",X"42",X"42",X"14",X"21",
		X"FC",X"00",X"08",X"00",X"08",X"00",X"04",X"00",X"01",X"F6",X"42",X"42",X"14",X"21",X"FE",X"00",
		X"FF",X"00",X"FF",X"00",X"C0",X"00",X"01",X"F6",X"42",X"42",X"14",X"21",X"FA",X"00",X"FF",X"00",
		X"E0",X"00",X"80",X"00",X"01",X"F6",X"42",X"42",X"14",X"21",X"F8",X"00",X"E0",X"00",X"C0",X"00",
		X"40",X"00",X"01",X"F6",X"42",X"42",X"14",X"21",X"F6",X"00",X"39",X"00",X"26",X"00",X"13",X"00",
		X"0C",X"F6",X"42",X"42",X"14",X"21",X"FE",X"00",X"2C",X"00",X"1C",X"00",X"0C",X"00",X"09",X"F6",
		X"42",X"42",X"14",X"21",X"FE",X"00",X"1F",X"00",X"13",X"00",X"09",X"00",X"06",X"F6",X"42",X"42",
		X"14",X"21",X"FC",X"00",X"18",X"00",X"10",X"00",X"08",X"00",X"04",X"FE",X"A6",X"A6",X"2A",X"62",
		X"FE",X"00",X"70",X"00",X"50",X"00",X"30",X"00",X"18",X"F6",X"42",X"42",X"14",X"21",X"FE",X"00",
		X"10",X"00",X"08",X"00",X"04",X"00",X"02",X"F6",X"42",X"42",X"14",X"21",X"FE",X"00",X"08",X"00",
		X"08",X"00",X"07",X"00",X"05",X"F6",X"42",X"42",X"14",X"21",X"FC",X"00",X"04",X"00",X"03",X"00",
		X"02",X"00",X"01",X"F6",X"42",X"42",X"14",X"21",X"FC",X"0A",X"8C",X"0A",X"8C",X"05",X"46",X"03",
		X"84",X"F6",X"42",X"42",X"14",X"21",X"88",X"00",X"18",X"00",X"10",X"00",X"08",X"00",X"00",X"FE",
		X"A6",X"A6",X"2A",X"62",X"FC",X"00",X"01",X"00",X"02",X"00",X"04",X"00",X"10",X"F6",X"42",X"42",
		X"14",X"21",X"04",X"01",X"0E",X"00",X"D2",X"00",X"96",X"00",X"3C",X"F6",X"42",X"42",X"14",X"21",
		X"F8",X"0B",X"9A",X"0A",X"8C",X"07",X"08",X"01",X"C2",X"F6",X"42",X"42",X"14",X"21",X"E2",X"0B",
		X"9A",X"0A",X"8C",X"07",X"08",X"01",X"C2",X"F6",X"42",X"42",X"14",X"21",X"E2",X"0B",X"9A",X"0A",
		X"8C",X"07",X"08",X"01",X"C2",X"F6",X"42",X"42",X"14",X"21",X"E2",X"00",X"30",X"00",X"28",X"00",
		X"20",X"00",X"10",X"F8",X"44",X"84",X"44",X"21",X"FC",X"00",X"02",X"00",X"02",X"00",X"03",X"00",
		X"0D",X"83",X"21",X"32",X"13",X"21",X"01",X"00",X"01",X"00",X"02",X"00",X"03",X"00",X"0D",X"95",
		X"32",X"53",X"25",X"32",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"0D",X"A7",X"53",X"75",
		X"37",X"53",X"01",X"8E",X"CC",X"14",X"BD",X"00",X"24",X"A7",X"E2",X"8E",X"14",X"2D",X"10",X"8E",
		X"B8",X"3B",X"E6",X"22",X"27",X"04",X"6A",X"22",X"26",X"2A",X"E6",X"E4",X"CB",X"10",X"57",X"E6",
		X"85",X"25",X"04",X"54",X"54",X"54",X"54",X"C4",X"0F",X"E7",X"22",X"E6",X"0D",X"1D",X"2B",X"09",
		X"E3",X"A4",X"10",X"A3",X"06",X"2D",X"0B",X"20",X"07",X"E3",X"A4",X"10",X"A3",X"06",X"2E",X"02",
		X"EC",X"06",X"ED",X"A4",X"30",X"0E",X"31",X"23",X"8C",X"16",X"33",X"25",X"C5",X"35",X"82",X"8E",
		X"19",X"33",X"20",X"03",X"8E",X"18",X"EA",X"EC",X"E1",X"34",X"10",X"ED",X"C8",X"12",X"8E",X"19",
		X"7C",X"10",X"8E",X"D0",X"10",X"F6",X"9A",X"4E",X"C4",X"0F",X"58",X"58",X"58",X"3A",X"EC",X"81",
		X"ED",X"A1",X"10",X"8C",X"D0",X"18",X"25",X"F6",X"4F",X"5F",X"ED",X"A1",X"ED",X"A1",X"ED",X"A1",
		X"ED",X"A1",X"35",X"06",X"DD",X"6F",X"8E",X"91",X"02",X"86",X"01",X"C6",X"FF",X"BD",X"18",X"C6",
		X"E7",X"80",X"4C",X"26",X"F6",X"CC",X"01",X"02",X"FD",X"9A",X"46",X"86",X"FF",X"B7",X"9A",X"49",
		X"86",X"01",X"B7",X"9A",X"45",X"B7",X"9A",X"43",X"86",X"08",X"B7",X"9A",X"44",X"FC",X"9A",X"4A",
		X"81",X"48",X"22",X"03",X"40",X"8B",X"90",X"1F",X"89",X"3D",X"34",X"06",X"86",X"F8",X"B0",X"9A",
		X"4B",X"44",X"1F",X"89",X"3D",X"E3",X"E4",X"ED",X"E4",X"8E",X"00",X"7F",X"30",X"1F",X"1F",X"10",
		X"1F",X"98",X"3D",X"A3",X"E4",X"22",X"F5",X"1F",X"10",X"CB",X"01",X"F7",X"9A",X"42",X"96",X"68",
		X"2B",X"07",X"BD",X"E0",X"A4",X"10",X"25",X"10",X"2E",X"8E",X"91",X"02",X"F6",X"9A",X"45",X"3A",
		X"A6",X"84",X"BD",X"17",X"62",X"B6",X"9A",X"49",X"80",X"11",X"81",X"88",X"24",X"02",X"86",X"FF",
		X"B7",X"9A",X"49",X"B6",X"9A",X"45",X"BB",X"9A",X"43",X"B7",X"9A",X"45",X"B1",X"9A",X"42",X"22",
		X"1E",X"7A",X"9A",X"44",X"26",X"C8",X"86",X"07",X"B7",X"9A",X"44",X"7C",X"9A",X"43",X"FC",X"9A",
		X"46",X"81",X"01",X"22",X"02",X"4F",X"5F",X"C3",X"02",X"04",X"FD",X"9A",X"46",X"20",X"AF",X"6E",
		X"D8",X"12",X"C6",X"FF",X"FD",X"9A",X"4C",X"10",X"8E",X"C8",X"80",X"8E",X"1A",X"7C",X"B6",X"9A",
		X"4D",X"E6",X"86",X"B6",X"9A",X"45",X"3D",X"34",X"02",X"8E",X"1B",X"7C",X"B6",X"9A",X"4D",X"E6",
		X"86",X"B6",X"9A",X"45",X"3D",X"E6",X"E4",X"34",X"02",X"58",X"34",X"06",X"1A",X"F0",X"FC",X"9A",
		X"46",X"ED",X"26",X"ED",X"22",X"B6",X"9A",X"49",X"A7",X"21",X"FC",X"9A",X"4A",X"A0",X"E4",X"25",
		X"5C",X"EB",X"61",X"25",X"3E",X"C1",X"F4",X"22",X"3A",X"ED",X"24",X"C6",X"12",X"E7",X"A4",X"F6",
		X"9A",X"4B",X"E0",X"61",X"25",X"1E",X"ED",X"24",X"86",X"12",X"A7",X"A4",X"B6",X"9A",X"4A",X"AB",
		X"E4",X"25",X"60",X"81",X"8E",X"22",X"5C",X"ED",X"24",X"C6",X"12",X"E7",X"A4",X"F6",X"9A",X"4B",
		X"EB",X"61",X"20",X"49",X"FC",X"9A",X"4A",X"AB",X"E4",X"25",X"48",X"81",X"8E",X"22",X"44",X"EB",
		X"61",X"20",X"3A",X"F6",X"9A",X"4B",X"E0",X"61",X"25",X"39",X"ED",X"24",X"86",X"12",X"A7",X"A4",
		X"B6",X"9A",X"4A",X"AB",X"E4",X"25",X"2C",X"81",X"8E",X"22",X"28",X"20",X"20",X"FC",X"9A",X"4A",
		X"AB",X"E4",X"25",X"1F",X"81",X"8E",X"22",X"1B",X"E0",X"61",X"25",X"06",X"ED",X"24",X"C6",X"12",
		X"E7",X"A4",X"F6",X"9A",X"4B",X"EB",X"61",X"25",X"0A",X"C1",X"F4",X"22",X"06",X"ED",X"24",X"C6",
		X"12",X"E7",X"A4",X"EC",X"62",X"1E",X"89",X"58",X"ED",X"E4",X"FC",X"9A",X"4A",X"A0",X"E4",X"25",
		X"5C",X"EB",X"61",X"25",X"3E",X"C1",X"F4",X"22",X"3A",X"ED",X"24",X"C6",X"12",X"E7",X"A4",X"F6",
		X"9A",X"4B",X"E0",X"61",X"25",X"1E",X"ED",X"24",X"86",X"12",X"A7",X"A4",X"B6",X"9A",X"4A",X"AB",
		X"E4",X"25",X"60",X"81",X"8E",X"22",X"5C",X"ED",X"24",X"C6",X"12",X"E7",X"A4",X"F6",X"9A",X"4B",
		X"EB",X"61",X"20",X"49",X"FC",X"9A",X"4A",X"AB",X"E4",X"25",X"48",X"81",X"8E",X"22",X"44",X"EB",
		X"61",X"20",X"3A",X"F6",X"9A",X"4B",X"E0",X"61",X"25",X"39",X"ED",X"24",X"86",X"12",X"A7",X"A4",
		X"B6",X"9A",X"4A",X"AB",X"E4",X"25",X"2C",X"81",X"8E",X"22",X"28",X"20",X"20",X"FC",X"9A",X"4A",
		X"AB",X"E4",X"25",X"1F",X"81",X"8E",X"22",X"1B",X"E0",X"61",X"25",X"06",X"ED",X"24",X"C6",X"12",
		X"E7",X"A4",X"F6",X"9A",X"4B",X"EB",X"61",X"25",X"0A",X"C1",X"F4",X"22",X"06",X"ED",X"24",X"C6",
		X"12",X"E7",X"A4",X"1C",X"EF",X"35",X"16",X"F6",X"9A",X"4D",X"F0",X"9A",X"4C",X"25",X"06",X"F7",
		X"9A",X"4D",X"7E",X"17",X"6B",X"39",X"34",X"06",X"4F",X"6F",X"61",X"58",X"5C",X"20",X"07",X"6C",
		X"61",X"A0",X"E4",X"58",X"27",X"09",X"49",X"68",X"61",X"A1",X"E4",X"25",X"F6",X"20",X"F0",X"48",
		X"25",X"04",X"A1",X"E4",X"25",X"02",X"6C",X"61",X"35",X"86",X"BE",X"D0",X"10",X"FC",X"D0",X"12",
		X"FD",X"D0",X"10",X"FD",X"80",X"F0",X"FC",X"D0",X"14",X"FD",X"D0",X"12",X"FD",X"80",X"F2",X"FC",
		X"D0",X"16",X"FD",X"D0",X"14",X"FD",X"80",X"F4",X"FC",X"D0",X"18",X"FD",X"D0",X"16",X"FD",X"80",
		X"F6",X"FC",X"D0",X"1A",X"FD",X"D0",X"18",X"FD",X"80",X"F8",X"FC",X"D0",X"1C",X"FD",X"D0",X"1A",
		X"FD",X"80",X"FA",X"FC",X"D0",X"1E",X"FD",X"D0",X"1C",X"FD",X"80",X"FC",X"BF",X"D0",X"1E",X"BF",
		X"80",X"FE",X"39",X"BE",X"D0",X"1E",X"FC",X"D0",X"1C",X"FD",X"D0",X"1E",X"FD",X"80",X"FE",X"FC",
		X"D0",X"1A",X"FD",X"D0",X"1C",X"FD",X"80",X"FC",X"FC",X"D0",X"18",X"FD",X"D0",X"1A",X"FD",X"80",
		X"FA",X"FC",X"D0",X"16",X"FD",X"D0",X"18",X"FD",X"80",X"F8",X"FC",X"D0",X"14",X"FD",X"D0",X"16",
		X"FD",X"80",X"F6",X"FC",X"D0",X"12",X"FD",X"D0",X"14",X"FD",X"80",X"F4",X"FC",X"D0",X"10",X"FD",
		X"D0",X"12",X"FD",X"80",X"F2",X"BF",X"D0",X"10",X"BF",X"80",X"F0",X"39",X"00",X"00",X"0E",X"D1",
		X"EE",X"C1",X"0E",X"D1",X"00",X"00",X"BB",X"DA",X"FF",X"DF",X"BB",X"DA",X"00",X"00",X"F0",X"B0",
		X"F0",X"F0",X"F0",X"B0",X"00",X"00",X"F0",X"B0",X"F0",X"F0",X"F0",X"B0",X"00",X"00",X"0F",X"B0",
		X"0F",X"F0",X"0F",X"B0",X"00",X"00",X"0F",X"B0",X"0F",X"F0",X"0F",X"B0",X"00",X"00",X"FF",X"B0",
		X"FF",X"F0",X"FF",X"B0",X"00",X"00",X"FF",X"B0",X"FF",X"F0",X"FF",X"B0",X"00",X"00",X"00",X"BF",
		X"00",X"FF",X"00",X"BF",X"00",X"00",X"0F",X"BF",X"0F",X"FF",X"0F",X"BF",X"00",X"00",X"0F",X"BF",
		X"0F",X"FF",X"0F",X"BF",X"00",X"00",X"F0",X"BF",X"F0",X"FF",X"F0",X"BF",X"00",X"00",X"F0",X"BF",
		X"F0",X"FF",X"F0",X"BF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"F0",X"F0",X"FF",X"FF",X"00",X"00",X"00",X"00",X"F0",X"FF",X"62",X"63",X"63",X"64",
		X"65",X"66",X"66",X"67",X"68",X"68",X"69",X"6A",X"6B",X"6B",X"6C",X"6D",X"6D",X"6E",X"6F",X"70",
		X"70",X"71",X"72",X"72",X"73",X"74",X"74",X"75",X"76",X"77",X"77",X"78",X"79",X"79",X"7A",X"7B",
		X"7B",X"7C",X"7D",X"7D",X"7E",X"7F",X"7F",X"80",X"81",X"82",X"82",X"83",X"84",X"84",X"85",X"86",
		X"86",X"87",X"88",X"88",X"89",X"8A",X"8A",X"8B",X"8C",X"8C",X"8D",X"8E",X"8E",X"8F",X"8F",X"90",
		X"91",X"91",X"92",X"93",X"93",X"94",X"95",X"95",X"96",X"97",X"97",X"98",X"98",X"99",X"9A",X"9A",
		X"9B",X"9C",X"9C",X"9D",X"9D",X"9E",X"9F",X"9F",X"A0",X"A0",X"A1",X"A2",X"A2",X"A3",X"A4",X"A4",
		X"A5",X"A5",X"A6",X"A7",X"A7",X"A8",X"A8",X"A9",X"A9",X"AA",X"AB",X"AB",X"AC",X"AC",X"AD",X"AE",
		X"AE",X"AF",X"AF",X"B0",X"B0",X"B1",X"B2",X"B2",X"B3",X"B3",X"B4",X"B4",X"00",X"01",X"02",X"02",
		X"03",X"04",X"05",X"05",X"06",X"07",X"08",X"09",X"09",X"0A",X"0B",X"0C",X"0D",X"0D",X"0E",X"0F",
		X"10",X"10",X"11",X"12",X"13",X"14",X"14",X"15",X"16",X"17",X"18",X"18",X"19",X"1A",X"1B",X"1B",
		X"1C",X"1D",X"1E",X"1F",X"1F",X"20",X"21",X"22",X"22",X"23",X"24",X"25",X"26",X"26",X"27",X"28",
		X"29",X"29",X"2A",X"2B",X"2C",X"2D",X"2D",X"2E",X"2F",X"30",X"30",X"31",X"32",X"33",X"33",X"34",
		X"35",X"36",X"37",X"37",X"38",X"39",X"3A",X"3A",X"3B",X"3C",X"3D",X"3D",X"3E",X"3F",X"40",X"40",
		X"41",X"42",X"43",X"44",X"44",X"45",X"46",X"47",X"47",X"48",X"49",X"4A",X"4A",X"4B",X"4C",X"4D",
		X"4D",X"4E",X"4F",X"50",X"50",X"51",X"52",X"53",X"53",X"54",X"55",X"55",X"56",X"57",X"58",X"58",
		X"59",X"5A",X"5B",X"5B",X"5C",X"5D",X"5E",X"5E",X"5F",X"60",X"60",X"61",X"EB",X"EB",X"EB",X"EB",
		X"EA",X"EA",X"EA",X"E9",X"E9",X"E9",X"E8",X"E8",X"E8",X"E7",X"E7",X"E7",X"E6",X"E6",X"E6",X"E5",
		X"E5",X"E5",X"E4",X"E4",X"E4",X"E3",X"E3",X"E2",X"E2",X"E2",X"E1",X"E1",X"E1",X"E0",X"E0",X"E0",
		X"DF",X"DF",X"DE",X"DE",X"DE",X"DD",X"DD",X"DC",X"DC",X"DC",X"DB",X"DB",X"DA",X"DA",X"DA",X"D9",
		X"D9",X"D8",X"D8",X"D8",X"D7",X"D7",X"D6",X"D6",X"D5",X"D5",X"D5",X"D4",X"D4",X"D3",X"D3",X"D2",
		X"D2",X"D1",X"D1",X"D1",X"D0",X"D0",X"CF",X"CF",X"CE",X"CE",X"CD",X"CD",X"CC",X"CC",X"CB",X"CB",
		X"CB",X"CA",X"CA",X"C9",X"C9",X"C8",X"C8",X"C7",X"C7",X"C6",X"C6",X"C5",X"C5",X"C4",X"C4",X"C3",
		X"C3",X"C2",X"C2",X"C1",X"C1",X"C0",X"C0",X"BF",X"BF",X"BE",X"BE",X"BD",X"BC",X"BC",X"BB",X"BB",
		X"BA",X"BA",X"B9",X"B9",X"B8",X"B8",X"B7",X"B7",X"B6",X"B5",X"B5",X"B4",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F8",X"F8",X"F8",X"F8",X"F8",X"F7",X"F7",X"F7",X"F7",X"F7",
		X"F7",X"F6",X"F6",X"F6",X"F6",X"F5",X"F5",X"F5",X"F5",X"F5",X"F4",X"F4",X"F4",X"F4",X"F3",X"F3",
		X"F3",X"F3",X"F3",X"F2",X"F2",X"F2",X"F2",X"F1",X"F1",X"F1",X"F1",X"F0",X"F0",X"F0",X"EF",X"EF",
		X"EF",X"EF",X"EE",X"EE",X"EE",X"ED",X"ED",X"ED",X"ED",X"EC",X"EC",X"EC",X"8E",X"30",X"90",X"CC",
		X"00",X"11",X"7E",X"E0",X"10",X"CC",X"00",X"F0",X"BD",X"E0",X"66",X"CC",X"11",X"FF",X"BD",X"E0",
		X"66",X"10",X"8E",X"27",X"1E",X"86",X"48",X"5F",X"BD",X"E0",X"63",X"7E",X"11",X"9E",X"0F",X"6E",
		X"20",X"4E",X"0F",X"68",X"86",X"80",X"97",X"6E",X"86",X"2C",X"A7",X"48",X"8D",X"CE",X"86",X"01",
		X"BD",X"E0",X"7D",X"6A",X"48",X"26",X"F5",X"10",X"8E",X"27",X"1E",X"86",X"48",X"5F",X"BD",X"E0",
		X"63",X"7E",X"00",X"54",X"0F",X"6E",X"96",X"E4",X"27",X"08",X"8E",X"29",X"8D",X"BD",X"E0",X"75",
		X"20",X"18",X"8E",X"29",X"95",X"BD",X"E0",X"75",X"96",X"90",X"2F",X"0E",X"6F",X"48",X"BD",X"1B",
		X"FC",X"86",X"01",X"BD",X"E0",X"7D",X"6A",X"48",X"26",X"F4",X"BD",X"E0",X"AD",X"BD",X"11",X"9E",
		X"0F",X"28",X"0F",X"68",X"CC",X"00",X"00",X"BD",X"E0",X"66",X"BD",X"E0",X"AD",X"BD",X"11",X"32",
		X"8E",X"24",X"64",X"BD",X"E0",X"6F",X"86",X"04",X"BD",X"E0",X"7D",X"BD",X"00",X"21",X"86",X"31",
		X"A7",X"51",X"B6",X"CC",X"05",X"46",X"24",X"75",X"CC",X"03",X"84",X"ED",X"48",X"8E",X"24",X"54",
		X"BD",X"E0",X"6F",X"8E",X"28",X"CE",X"AF",X"4A",X"BD",X"28",X"94",X"86",X"02",X"BD",X"E0",X"7D",
		X"CE",X"29",X"32",X"10",X"8E",X"29",X"1E",X"AE",X"C4",X"E6",X"43",X"A6",X"42",X"BD",X"29",X"04",
		X"4A",X"26",X"FA",X"A6",X"21",X"34",X"02",X"1E",X"10",X"A6",X"C4",X"EB",X"E0",X"1E",X"01",X"5A",
		X"26",X"E9",X"33",X"44",X"11",X"83",X"29",X"5E",X"25",X"DD",X"BD",X"00",X"36",X"BD",X"25",X"59",
		X"86",X"01",X"BD",X"E0",X"7D",X"BD",X"28",X"94",X"7C",X"D0",X"04",X"EC",X"48",X"C3",X"FF",X"FF",
		X"ED",X"48",X"26",X"EC",X"BD",X"26",X"83",X"83",X"00",X"03",X"26",X"07",X"CC",X"00",X"3C",X"ED",
		X"48",X"20",X"DD",X"10",X"8E",X"24",X"44",X"86",X"49",X"5F",X"BD",X"E0",X"63",X"BD",X"E0",X"AA",
		X"BD",X"11",X"20",X"8E",X"24",X"A4",X"BD",X"E0",X"6F",X"86",X"02",X"BD",X"E0",X"7D",X"34",X"01",
		X"1A",X"F0",X"86",X"22",X"B7",X"C8",X"81",X"CC",X"90",X"01",X"FD",X"C8",X"86",X"CC",X"00",X"BA",
		X"FD",X"C8",X"84",X"86",X"12",X"B7",X"C8",X"80",X"C6",X"E1",X"F7",X"C8",X"85",X"B7",X"C8",X"80",
		X"35",X"01",X"BD",X"00",X"51",X"CC",X"19",X"1A",X"BD",X"1E",X"32",X"86",X"10",X"BD",X"E0",X"7D",
		X"CC",X"1B",X"1C",X"BD",X"1E",X"32",X"86",X"04",X"BD",X"E0",X"7D",X"CC",X"1D",X"1E",X"BD",X"1E",
		X"32",X"31",X"48",X"8E",X"1D",X"FB",X"A6",X"80",X"A7",X"A0",X"8C",X"1E",X"1E",X"25",X"F7",X"86",
		X"01",X"BD",X"E0",X"7D",X"C6",X"07",X"33",X"48",X"A6",X"44",X"2B",X"1C",X"26",X"18",X"AE",X"C4",
		X"10",X"AE",X"42",X"34",X"04",X"86",X"02",X"BD",X"E0",X"99",X"38",X"00",X"05",X"35",X"04",X"AF",
		X"C4",X"10",X"AF",X"42",X"24",X"02",X"6A",X"44",X"33",X"45",X"5A",X"26",X"DB",X"A6",X"5F",X"2A",
		X"CE",X"CC",X"C0",X"51",X"FD",X"B8",X"18",X"86",X"0F",X"B7",X"B8",X"23",X"10",X"8E",X"30",X"26",
		X"CC",X"0F",X"FF",X"BD",X"E0",X"63",X"8E",X"00",X"BC",X"CC",X"58",X"77",X"BD",X"E0",X"56",X"10",
		X"8E",X"1E",X"1E",X"86",X"90",X"5F",X"BD",X"E0",X"63",X"86",X"F0",X"BD",X"E0",X"7D",X"86",X"F0",
		X"BD",X"E0",X"7D",X"86",X"F0",X"BD",X"E0",X"7D",X"CC",X"47",X"20",X"FD",X"9A",X"4A",X"BD",X"E0",
		X"72",X"B7",X"9A",X"4E",X"CC",X"90",X"FF",X"BD",X"E0",X"66",X"CC",X"0F",X"FF",X"BD",X"E0",X"66",
		X"BD",X"16",X"84",X"86",X"3C",X"BD",X"E0",X"7D",X"7E",X"1E",X"3D",X"55",X"28",X"38",X"03",X"02",
		X"5A",X"28",X"39",X"66",X"0C",X"66",X"28",X"3C",X"44",X"16",X"73",X"28",X"3E",X"04",X"20",X"80",
		X"28",X"3F",X"B4",X"2A",X"8D",X"28",X"42",X"B4",X"34",X"9F",X"28",X"45",X"E9",X"3E",X"BD",X"E0",
		X"99",X"EF",X"E0",X"05",X"BD",X"E0",X"99",X"EF",X"E3",X"05",X"8E",X"1E",X"24",X"86",X"01",X"7E",
		X"E0",X"6C",X"FD",X"C0",X"51",X"88",X"80",X"C8",X"80",X"FD",X"C0",X"61",X"39",X"7F",X"B8",X"AA",
		X"86",X"7F",X"97",X"68",X"86",X"05",X"97",X"4A",X"97",X"49",X"7E",X"27",X"C1",X"10",X"8E",X"24",
		X"44",X"86",X"49",X"5F",X"BD",X"E0",X"63",X"4F",X"5F",X"DD",X"69",X"BD",X"25",X"59",X"8E",X"1E",
		X"F4",X"AF",X"48",X"6F",X"4B",X"6F",X"4D",X"6F",X"4F",X"6F",X"C8",X"11",X"6F",X"C8",X"13",X"AE",
		X"48",X"30",X"06",X"AF",X"48",X"8C",X"20",X"0E",X"10",X"24",X"FD",X"F4",X"A6",X"04",X"27",X"19",
		X"31",X"4B",X"8E",X"00",X"90",X"30",X"88",X"10",X"A1",X"A1",X"26",X"F9",X"5F",X"6F",X"3E",X"BD",
		X"E0",X"56",X"30",X"88",X"10",X"A6",X"A1",X"26",X"F3",X"86",X"02",X"BD",X"E0",X"7D",X"AE",X"48",
		X"A6",X"02",X"27",X"13",X"E6",X"03",X"31",X"4B",X"8E",X"00",X"90",X"30",X"88",X"10",X"6D",X"A1",
		X"26",X"F9",X"ED",X"3E",X"BD",X"E0",X"56",X"86",X"02",X"BD",X"E0",X"7D",X"AE",X"48",X"AD",X"94",
		X"AE",X"48",X"A6",X"05",X"27",X"A9",X"A7",X"4A",X"86",X"01",X"8D",X"12",X"86",X"02",X"8D",X"0E",
		X"86",X"03",X"8D",X"0A",X"86",X"04",X"8D",X"06",X"6A",X"4A",X"26",X"EC",X"20",X"91",X"31",X"49",
		X"8E",X"00",X"90",X"30",X"88",X"10",X"31",X"22",X"4A",X"26",X"F8",X"A6",X"A4",X"27",X"05",X"E6",
		X"21",X"BD",X"E0",X"56",X"86",X"04",X"7E",X"E0",X"7D",X"39",X"1E",X"F9",X"72",X"55",X"00",X"03",
		X"1E",X"F9",X"73",X"55",X"00",X"03",X"1E",X"F9",X"74",X"55",X"00",X"0A",X"20",X"0E",X"75",X"55",
		X"72",X"05",X"20",X"37",X"76",X"55",X"00",X"05",X"20",X"B2",X"77",X"55",X"00",X"05",X"20",X"7D",
		X"78",X"55",X"00",X"0A",X"20",X"E3",X"79",X"55",X"75",X"03",X"1E",X"F9",X"7A",X"55",X"00",X"03",
		X"1E",X"F9",X"7B",X"55",X"00",X"03",X"1E",X"F9",X"7C",X"55",X"00",X"0A",X"1E",X"F9",X"7D",X"55",
		X"79",X"03",X"1E",X"F9",X"7E",X"55",X"00",X"03",X"1E",X"F9",X"7F",X"55",X"00",X"0A",X"21",X"C7",
		X"80",X"55",X"7D",X"03",X"1E",X"F9",X"81",X"55",X"00",X"03",X"1E",X"F9",X"82",X"55",X"00",X"0A",
		X"22",X"61",X"83",X"33",X"80",X"01",X"22",X"6A",X"00",X"33",X"00",X"01",X"22",X"73",X"00",X"33",
		X"00",X"01",X"1E",X"F9",X"84",X"33",X"00",X"03",X"22",X"7C",X"85",X"CC",X"00",X"06",X"22",X"84",
		X"86",X"AA",X"85",X"06",X"22",X"91",X"87",X"EE",X"86",X"01",X"22",X"B3",X"00",X"EE",X"00",X"01",
		X"22",X"BC",X"00",X"EE",X"00",X"04",X"22",X"C8",X"88",X"33",X"83",X"03",X"23",X"11",X"89",X"33",
		X"00",X"03",X"23",X"07",X"8A",X"33",X"00",X"03",X"1E",X"F9",X"AB",X"99",X"00",X"0A",X"23",X"28",
		X"90",X"11",X"88",X"03",X"1E",X"F9",X"91",X"55",X"00",X"03",X"1E",X"F9",X"92",X"55",X"00",X"03",
		X"1E",X"F9",X"9D",X"55",X"00",X"0A",X"23",X"4B",X"93",X"BB",X"90",X"03",X"1E",X"F9",X"94",X"BB",
		X"00",X"03",X"23",X"59",X"95",X"BB",X"00",X"02",X"23",X"77",X"00",X"BB",X"00",X"01",X"1E",X"F9",
		X"96",X"BB",X"00",X"0A",X"23",X"C1",X"97",X"77",X"93",X"03",X"1E",X"F9",X"98",X"77",X"00",X"03",
		X"1E",X"F9",X"99",X"77",X"00",X"0A",X"23",X"E6",X"9A",X"EE",X"97",X"03",X"1E",X"F9",X"9B",X"EE",
		X"00",X"03",X"1E",X"F9",X"9C",X"EE",X"00",X"0A",X"23",X"EC",X"00",X"EE",X"9A",X"0A",X"BD",X"24",
		X"34",X"CC",X"21",X"8C",X"ED",X"A8",X"25",X"6F",X"A8",X"33",X"CC",X"20",X"21",X"ED",X"A8",X"37",
		X"39",X"01",X"19",X"1D",X"01",X"19",X"1F",X"01",X"17",X"1F",X"01",X"17",X"1B",X"01",X"15",X"1B",
		X"01",X"15",X"1D",X"01",X"17",X"1D",X"FF",X"BD",X"24",X"34",X"CC",X"20",X"4D",X"ED",X"A8",X"25",
		X"6F",X"23",X"CC",X"20",X"4E",X"ED",X"A8",X"27",X"4F",X"5F",X"ED",X"A8",X"33",X"39",X"6A",X"C8",
		X"33",X"2E",X"1B",X"8E",X"20",X"6F",X"E6",X"C8",X"34",X"3A",X"3A",X"6C",X"C8",X"34",X"EC",X"84",
		X"E7",X"C8",X"33",X"26",X"06",X"8E",X"20",X"4D",X"AF",X"C8",X"27",X"A7",X"C8",X"21",X"39",X"01",
		X"0A",X"02",X"05",X"08",X"08",X"02",X"05",X"01",X"08",X"02",X"7F",X"00",X"00",X"BD",X"24",X"34",
		X"CC",X"20",X"8A",X"ED",X"A8",X"27",X"6F",X"A8",X"39",X"39",X"6A",X"C8",X"39",X"2E",X"14",X"86",
		X"0C",X"A7",X"C8",X"39",X"A6",X"C8",X"10",X"8E",X"20",X"A9",X"E6",X"86",X"E7",X"C8",X"21",X"6C",
		X"C8",X"12",X"39",X"6F",X"C8",X"12",X"6F",X"C8",X"21",X"39",X"04",X"01",X"00",X"08",X"00",X"00",
		X"00",X"02",X"BD",X"24",X"34",X"CC",X"20",X"C7",X"ED",X"A8",X"27",X"C6",X"03",X"E7",X"A8",X"33",
		X"CC",X"20",X"C6",X"ED",X"A8",X"25",X"39",X"A6",X"C8",X"3B",X"26",X"10",X"6A",X"C8",X"33",X"26",
		X"07",X"CC",X"20",X"D7",X"ED",X"C8",X"27",X"39",X"6C",X"C8",X"12",X"39",X"6F",X"C8",X"12",X"6F",
		X"C8",X"21",X"39",X"BD",X"24",X"34",X"86",X"01",X"A7",X"A8",X"12",X"CC",X"21",X"01",X"ED",X"A8",
		X"27",X"CC",X"21",X"8C",X"ED",X"A8",X"25",X"6F",X"A8",X"33",X"CC",X"21",X"2B",X"ED",X"A8",X"37",
		X"39",X"FC",X"B7",X"18",X"2B",X"24",X"6F",X"C8",X"12",X"CC",X"21",X"10",X"ED",X"C8",X"27",X"39",
		X"10",X"BE",X"B7",X"18",X"2A",X"14",X"CC",X"21",X"32",X"ED",X"A8",X"27",X"86",X"08",X"A7",X"A8",
		X"21",X"6C",X"A8",X"12",X"CC",X"21",X"2A",X"ED",X"C8",X"27",X"39",X"01",X"1D",X"1D",X"01",X"1D",
		X"1B",X"FF",X"BE",X"B7",X"16",X"2B",X"F3",X"86",X"08",X"A7",X"43",X"EC",X"C8",X"16",X"83",X"1D",
		X"15",X"27",X"E7",X"86",X"02",X"A7",X"C8",X"21",X"CC",X"21",X"62",X"ED",X"C8",X"27",X"CC",X"21",
		X"8C",X"ED",X"C8",X"25",X"6F",X"C8",X"33",X"CC",X"21",X"85",X"ED",X"C8",X"37",X"86",X"1F",X"A7",
		X"C8",X"39",X"A6",X"C8",X"12",X"26",X"1A",X"A6",X"C8",X"3B",X"26",X"BE",X"6A",X"C8",X"39",X"26",
		X"0C",X"CC",X"21",X"2A",X"6F",X"43",X"ED",X"C8",X"25",X"ED",X"C8",X"27",X"39",X"6C",X"C8",X"12",
		X"39",X"6F",X"C8",X"12",X"39",X"08",X"1D",X"1D",X"02",X"1B",X"1D",X"FF",X"E6",X"C8",X"33",X"26",
		X"15",X"AE",X"C8",X"37",X"A6",X"80",X"2B",X"2C",X"A7",X"C8",X"21",X"EC",X"81",X"ED",X"C8",X"33",
		X"AF",X"C8",X"37",X"E6",X"C8",X"33",X"86",X"02",X"E0",X"C8",X"16",X"26",X"11",X"86",X"01",X"E6",
		X"C8",X"34",X"E0",X"C8",X"17",X"27",X"DA",X"2B",X"02",X"86",X"08",X"A7",X"43",X"39",X"2B",X"FB",
		X"86",X"04",X"20",X"F7",X"6F",X"43",X"39",X"BD",X"24",X"3C",X"CC",X"21",X"F1",X"ED",X"A8",X"25",
		X"6F",X"A8",X"33",X"CC",X"22",X"4F",X"ED",X"A8",X"37",X"BD",X"24",X"34",X"CC",X"22",X"25",X"ED",
		X"A8",X"25",X"6F",X"A8",X"33",X"CC",X"22",X"5D",X"ED",X"A8",X"37",X"86",X"05",X"A7",X"A8",X"39",
		X"39",X"FC",X"22",X"53",X"A3",X"C8",X"16",X"27",X"03",X"7E",X"21",X"8C",X"6F",X"43",X"6F",X"C8",
		X"21",X"A6",X"C8",X"12",X"27",X"48",X"CC",X"22",X"0D",X"ED",X"C8",X"25",X"39",X"6F",X"C8",X"12",
		X"A6",X"C8",X"3B",X"26",X"39",X"CC",X"22",X"56",X"ED",X"C8",X"37",X"6F",X"C8",X"33",X"CC",X"21",
		X"8C",X"ED",X"C8",X"25",X"39",X"FC",X"22",X"5E",X"A3",X"C8",X"16",X"27",X"03",X"7E",X"21",X"8C",
		X"6F",X"43",X"A6",X"C8",X"12",X"26",X"14",X"A6",X"C8",X"3B",X"26",X"12",X"6A",X"C8",X"39",X"26",
		X"06",X"BD",X"24",X"3C",X"6C",X"A8",X"12",X"6C",X"C8",X"12",X"39",X"6F",X"C8",X"12",X"39",X"02",
		X"1B",X"1D",X"02",X"16",X"1D",X"FF",X"02",X"1D",X"1D",X"01",X"1D",X"15",X"FF",X"04",X"11",X"1D",
		X"FF",X"7A",X"B7",X"73",X"86",X"0F",X"B7",X"B8",X"23",X"39",X"CC",X"1B",X"9B",X"8E",X"1C",X"9C",
		X"7E",X"30",X"20",X"CC",X"1D",X"9D",X"8E",X"1E",X"9E",X"7E",X"30",X"20",X"BD",X"30",X"0E",X"CC",
		X"04",X"62",X"20",X"06",X"BD",X"30",X"11",X"CC",X"04",X"5E",X"B3",X"91",X"00",X"ED",X"A8",X"41",
		X"39",X"BD",X"30",X"14",X"CC",X"04",X"5A",X"8D",X"F1",X"BD",X"24",X"34",X"CC",X"21",X"8C",X"ED",
		X"A8",X"25",X"CC",X"22",X"AC",X"ED",X"A8",X"37",X"6F",X"A8",X"33",X"39",X"02",X"13",X"1D",X"01",
		X"11",X"1D",X"FF",X"CC",X"1B",X"9B",X"8E",X"1C",X"9C",X"7E",X"30",X"20",X"7F",X"B8",X"23",X"CC",
		X"19",X"99",X"8E",X"1A",X"9A",X"7E",X"30",X"20",X"BD",X"24",X"34",X"CC",X"22",X"D2",X"ED",X"A8",
		X"25",X"39",X"A6",X"43",X"10",X"26",X"FE",X"B4",X"86",X"01",X"A7",X"C8",X"12",X"CC",X"22",X"E4",
		X"ED",X"C8",X"25",X"39",X"6F",X"C8",X"12",X"A6",X"C8",X"3B",X"26",X"1A",X"86",X"08",X"A7",X"C8",
		X"21",X"86",X"01",X"A7",X"C8",X"12",X"CC",X"22",X"FD",X"ED",X"C8",X"25",X"39",X"6F",X"C8",X"12",
		X"CC",X"23",X"06",X"ED",X"C8",X"25",X"39",X"BE",X"B7",X"1E",X"CC",X"30",X"23",X"ED",X"88",X"25",
		X"39",X"BD",X"24",X"34",X"CC",X"21",X"8C",X"ED",X"A8",X"25",X"CC",X"23",X"24",X"ED",X"A8",X"37",
		X"6F",X"A8",X"33",X"39",X"08",X"11",X"23",X"FF",X"BD",X"24",X"34",X"CC",X"23",X"35",X"ED",X"A8",
		X"37",X"6F",X"A8",X"33",X"39",X"02",X"0F",X"23",X"04",X"11",X"23",X"01",X"11",X"21",X"04",X"13",
		X"21",X"02",X"13",X"1F",X"02",X"15",X"1F",X"02",X"15",X"1D",X"FF",X"10",X"8E",X"30",X"17",X"86",
		X"04",X"C6",X"FF",X"BD",X"E0",X"63",X"0C",X"90",X"39",X"BD",X"24",X"34",X"CC",X"23",X"63",X"ED",
		X"A8",X"25",X"39",X"6F",X"C8",X"12",X"10",X"BE",X"B7",X"34",X"2A",X"0A",X"EC",X"A8",X"16",X"81",
		X"11",X"25",X"03",X"6C",X"C8",X"12",X"39",X"10",X"BE",X"B7",X"34",X"A6",X"A8",X"51",X"81",X"03",
		X"26",X"07",X"AE",X"48",X"30",X"1A",X"AF",X"48",X"39",X"BD",X"24",X"34",X"CC",X"23",X"9C",X"ED",
		X"A8",X"25",X"CC",X"23",X"B4",X"ED",X"A8",X"37",X"6F",X"A8",X"33",X"39",X"FC",X"23",X"BE",X"10",
		X"A3",X"C8",X"16",X"27",X"03",X"7E",X"21",X"8C",X"6F",X"43",X"10",X"BE",X"B7",X"34",X"2B",X"03",
		X"6F",X"C8",X"12",X"39",X"08",X"13",X"1D",X"08",X"13",X"19",X"08",X"11",X"19",X"08",X"11",X"1C",
		X"FF",X"10",X"BE",X"B7",X"34",X"10",X"2B",X"F8",X"A7",X"BD",X"24",X"34",X"CC",X"21",X"8C",X"ED",
		X"A8",X"25",X"CC",X"23",X"DC",X"ED",X"A8",X"37",X"6F",X"A8",X"33",X"39",X"08",X"11",X"1D",X"02",
		X"0D",X"1D",X"02",X"1D",X"0D",X"FF",X"7F",X"B7",X"73",X"7E",X"30",X"1A",X"10",X"8E",X"23",X"F7",
		X"86",X"60",X"5F",X"BD",X"E0",X"63",X"39",X"86",X"1E",X"BD",X"E0",X"7D",X"8E",X"CC",X"00",X"BD",
		X"00",X"24",X"4D",X"27",X"2C",X"CC",X"2D",X"55",X"8E",X"26",X"D0",X"BD",X"E0",X"10",X"34",X"10",
		X"8E",X"CC",X"00",X"BD",X"00",X"24",X"35",X"10",X"85",X"F0",X"26",X"06",X"8A",X"F0",X"30",X"89",
		X"FD",X"00",X"BD",X"E0",X"17",X"86",X"A0",X"BD",X"E0",X"10",X"86",X"04",X"BD",X"E0",X"7D",X"20",
		X"D4",X"7E",X"E0",X"69",X"10",X"BE",X"B7",X"16",X"2B",X"01",X"3F",X"39",X"10",X"BE",X"B7",X"18",
		X"2B",X"01",X"3F",X"39",X"86",X"05",X"BD",X"E0",X"7D",X"BD",X"26",X"83",X"83",X"00",X"03",X"26",
		X"F3",X"7E",X"1C",X"70",X"00",X"00",X"F0",X"B0",X"00",X"BF",X"0C",X"C7",X"00",X"BF",X"AE",X"D1",
		X"BB",X"DA",X"A0",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AE",X"D1",X"0F",X"90",X"0F",X"40",X"00",X"BF",X"AE",X"D1",
		X"BB",X"DA",X"A0",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"AF",X"BC",X"AC",X"B1",X"9A",X"BC",X"8B",X"BC",X"7B",
		X"BC",X"6B",X"CF",X"39",X"CF",X"59",X"CF",X"49",X"DF",X"2E",X"CD",X"7B",X"FF",X"8B",X"CC",X"AC",
		X"CC",X"9C",X"CC",X"8C",X"86",X"04",X"BD",X"E0",X"7D",X"86",X"1E",X"A7",X"48",X"BD",X"11",X"9E",
		X"8E",X"25",X"11",X"BD",X"E0",X"6F",X"BD",X"25",X"59",X"86",X"11",X"D6",X"E1",X"5A",X"27",X"02",
		X"86",X"12",X"BD",X"E0",X"33",X"86",X"3C",X"BD",X"E0",X"7D",X"6A",X"48",X"26",X"F7",X"7E",X"1C",
		X"70",X"00",X"00",X"FF",X"DF",X"75",X"CE",X"85",X"AE",X"A2",X"6F",X"AE",X"D1",X"BB",X"DA",X"EE",
		X"C1",X"00",X"00",X"0E",X"D1",X"0F",X"90",X"C0",X"D0",X"D8",X"A9",X"E2",X"50",X"6A",X"DA",X"19",
		X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"8E",X"29",X"92",X"BD",X"E0",X"75",X"0C",X"6E",X"8D",X"14",X"CC",X"4D",X"22",X"8E",X"38",
		X"E3",X"BD",X"E0",X"10",X"96",X"E1",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"7E",X"E0",X"17",X"34",
		X"01",X"1A",X"F0",X"CC",X"1F",X"09",X"FD",X"C8",X"86",X"CC",X"37",X"E2",X"FD",X"C8",X"84",X"FD",
		X"C8",X"82",X"7F",X"C8",X"81",X"86",X"12",X"B7",X"C8",X"80",X"35",X"81",X"34",X"76",X"CE",X"90",
		X"02",X"10",X"8E",X"25",X"9D",X"86",X"80",X"5F",X"BD",X"E0",X"78",X"35",X"F6",X"CC",X"80",X"FF",
		X"BD",X"E0",X"66",X"86",X"F0",X"D6",X"28",X"27",X"01",X"44",X"A7",X"48",X"8D",X"AB",X"86",X"01",
		X"BD",X"E0",X"7D",X"8D",X"A6",X"6A",X"48",X"26",X"F5",X"86",X"01",X"BD",X"E0",X"7D",X"CC",X"4D",
		X"00",X"8D",X"9B",X"7E",X"E0",X"69",X"96",X"6D",X"81",X"02",X"25",X"03",X"7E",X"E0",X"69",X"86",
		X"1E",X"BD",X"E0",X"7D",X"CC",X"00",X"C3",X"BD",X"26",X"6D",X"26",X"EA",X"BD",X"26",X"6D",X"27",
		X"FB",X"86",X"0F",X"BD",X"E0",X"7D",X"CC",X"00",X"C0",X"BD",X"26",X"6D",X"26",X"D8",X"BD",X"26",
		X"6D",X"27",X"FB",X"86",X"0F",X"BD",X"E0",X"7D",X"CC",X"00",X"41",X"BD",X"26",X"6D",X"26",X"C6",
		X"BD",X"26",X"6D",X"27",X"FB",X"86",X"0F",X"BD",X"E0",X"7D",X"CC",X"00",X"03",X"BD",X"26",X"6D",
		X"26",X"B4",X"BD",X"E0",X"AA",X"BD",X"00",X"21",X"1A",X"FF",X"86",X"03",X"B7",X"BF",X"FF",X"B7",
		X"C8",X"00",X"4F",X"5F",X"FD",X"80",X"00",X"4A",X"5A",X"FD",X"80",X"02",X"86",X"01",X"B7",X"BF",
		X"FF",X"B7",X"C8",X"00",X"CE",X"26",X"B0",X"8E",X"10",X"30",X"34",X"10",X"C6",X"11",X"A6",X"C0",
		X"88",X"9B",X"80",X"35",X"2B",X"10",X"27",X"05",X"BD",X"E0",X"09",X"20",X"F1",X"AE",X"E4",X"30",
		X"88",X"10",X"AF",X"E4",X"20",X"E8",X"8E",X"1B",X"E6",X"86",X"14",X"B7",X"C9",X"00",X"8D",X"23",
		X"83",X"00",X"03",X"27",X"F1",X"30",X"1F",X"26",X"F0",X"6E",X"9F",X"EF",X"FE",X"ED",X"48",X"EC",
		X"E1",X"ED",X"4A",X"86",X"01",X"BD",X"E0",X"7D",X"8D",X"09",X"1F",X"01",X"EC",X"48",X"AC",X"48",
		X"6E",X"D8",X"0A",X"F6",X"C9",X"86",X"C4",X"C0",X"B6",X"C9",X"85",X"84",X"C7",X"8A",X"30",X"B7",
		X"C9",X"85",X"B6",X"C9",X"84",X"43",X"84",X"30",X"27",X"02",X"CA",X"01",X"B6",X"C9",X"85",X"8A",
		X"38",X"B7",X"C9",X"85",X"B6",X"C9",X"84",X"43",X"84",X"30",X"27",X"02",X"CA",X"02",X"4F",X"39",
		X"C8",X"DC",X"D3",X"C9",X"A4",X"D3",X"C9",X"A4",X"D3",X"D6",X"DE",X"DF",X"CA",X"D6",X"D5",X"AE",
		X"D8",X"DF",X"C9",X"D3",X"DD",X"D6",X"DF",X"D8",X"A4",X"DA",X"C3",X"A4",X"CD",X"D3",X"D0",X"D0",
		X"D3",X"DB",X"D7",X"C9",X"A4",X"DF",X"D0",X"DF",X"D9",X"C8",X"CA",X"D5",X"D6",X"D3",X"D9",X"C9",
		X"A4",X"D3",X"D6",X"D9",X"F8",X"AE",X"C4",X"D9",X"FB",X"A4",X"AD",X"A5",X"A6",X"A2",X"A4",X"CD",
		X"D3",X"D0",X"D0",X"D3",X"DB",X"D7",X"C9",X"A4",X"DF",X"D0",X"DF",X"D9",X"C8",X"CA",X"D5",X"D6",
		X"D3",X"D9",X"C9",X"A4",X"D3",X"D6",X"D9",X"F8",X"AE",X"DB",X"D0",X"D0",X"A4",X"CA",X"D3",X"DD",
		X"DC",X"C8",X"C9",X"A4",X"CA",X"DF",X"C9",X"DF",X"CA",X"CE",X"DF",X"CA",X"D8",X"2E",X"CC",X"48",
		X"FF",X"BD",X"E0",X"66",X"86",X"01",X"BD",X"E0",X"7D",X"96",X"6E",X"2F",X"15",X"0F",X"6E",X"CC",
		X"00",X"00",X"BD",X"E0",X"66",X"BD",X"E0",X"AD",X"10",X"8E",X"24",X"E4",X"86",X"47",X"5F",X"BD",
		X"E0",X"63",X"BD",X"E0",X"A4",X"24",X"DD",X"8E",X"CC",X"06",X"BD",X"00",X"24",X"81",X"09",X"27",
		X"10",X"1F",X"98",X"40",X"8B",X"99",X"9B",X"E1",X"19",X"97",X"E1",X"8E",X"CD",X"00",X"BD",X"00",
		X"2D",X"86",X"08",X"0F",X"49",X"5D",X"27",X"09",X"86",X"09",X"0C",X"49",X"C6",X"0B",X"BD",X"00",
		X"1E",X"1F",X"89",X"BD",X"00",X"1E",X"C6",X"0B",X"BD",X"00",X"1E",X"C6",X"07",X"BD",X"00",X"1E",
		X"7F",X"B8",X"AA",X"8E",X"CC",X"02",X"BD",X"00",X"27",X"D7",X"4A",X"CC",X"00",X"00",X"BD",X"E0",
		X"66",X"BD",X"E0",X"AD",X"0F",X"4C",X"86",X"FF",X"97",X"68",X"8E",X"29",X"8A",X"BD",X"E0",X"75",
		X"CC",X"91",X"BD",X"83",X"68",X"23",X"1F",X"01",X"CC",X"00",X"2C",X"AB",X"80",X"5A",X"26",X"FB",
		X"80",X"00",X"27",X"03",X"7C",X"B8",X"AA",X"10",X"8E",X"25",X"C6",X"86",X"50",X"5F",X"BD",X"E0",
		X"63",X"86",X"04",X"BD",X"E0",X"7D",X"BD",X"E0",X"AA",X"BD",X"00",X"21",X"0F",X"6D",X"BE",X"E0",
		X"7B",X"BD",X"E0",X"6F",X"CE",X"28",X"73",X"AE",X"C1",X"EC",X"C1",X"80",X"21",X"88",X"12",X"BD",
		X"E0",X"09",X"A6",X"C0",X"26",X"F5",X"DE",X"21",X"8E",X"90",X"2B",X"6F",X"80",X"8C",X"90",X"49",
		X"25",X"F9",X"8E",X"CC",X"00",X"BD",X"00",X"27",X"4F",X"58",X"49",X"58",X"49",X"58",X"49",X"58",
		X"49",X"DD",X"69",X"DD",X"34",X"DD",X"43",X"8E",X"CC",X"14",X"BD",X"00",X"24",X"6F",X"E2",X"81",
		X"03",X"23",X"08",X"6C",X"E4",X"81",X"06",X"23",X"02",X"6C",X"E4",X"8E",X"14",X"2D",X"10",X"8E",
		X"B8",X"3B",X"E6",X"E4",X"58",X"EC",X"85",X"ED",X"A4",X"86",X"02",X"A7",X"22",X"30",X"0E",X"31",
		X"23",X"8C",X"16",X"33",X"25",X"EC",X"D6",X"4A",X"BD",X"00",X"48",X"96",X"4A",X"8B",X"99",X"19",
		X"97",X"30",X"D7",X"31",X"0D",X"49",X"27",X"04",X"97",X"3F",X"D7",X"40",X"10",X"8E",X"13",X"08",
		X"86",X"21",X"C6",X"FF",X"BD",X"E0",X"63",X"CC",X"12",X"8C",X"ED",X"28",X"96",X"49",X"27",X"10",
		X"10",X"8E",X"13",X"08",X"86",X"22",X"C6",X"FF",X"BD",X"E0",X"63",X"CC",X"12",X"CA",X"ED",X"28",
		X"7E",X"30",X"00",X"10",X"F8",X"59",X"11",X"40",X"5A",X"39",X"54",X"22",X"25",X"25",X"22",X"3A",
		X"26",X"30",X"39",X"3E",X"25",X"3E",X"40",X"2D",X"2F",X"2C",X"2B",X"22",X"40",X"30",X"39",X"22",
		X"2B",X"40",X"5D",X"00",X"AE",X"4A",X"EC",X"81",X"FD",X"D0",X"1E",X"EC",X"81",X"FD",X"D0",X"1C",
		X"EC",X"81",X"FD",X"D0",X"1A",X"EC",X"81",X"FD",X"D0",X"18",X"EC",X"81",X"FD",X"D0",X"16",X"EC",
		X"81",X"FD",X"D0",X"14",X"EC",X"81",X"FD",X"D0",X"12",X"EC",X"81",X"FD",X"D0",X"10",X"EC",X"81",
		X"FD",X"D0",X"0E",X"8C",X"29",X"04",X"25",X"03",X"8E",X"28",X"CE",X"AF",X"4A",X"39",X"00",X"DF",
		X"00",X"DF",X"00",X"00",X"00",X"DF",X"00",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"DF",X"00",X"DF",X"00",X"00",X"00",X"DF",X"00",X"DF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"DF",X"00",X"00",X"00",X"DF",X"00",X"DF",X"00",X"00",X"00",X"DF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"34",X"27",X"1A",X"F0",X"EC",X"A1",X"FD",X"C8",X"86",X"BF",X"C8",X"84",
		X"10",X"BF",X"C8",X"82",X"C6",X"02",X"F7",X"C8",X"80",X"5F",X"30",X"8B",X"35",X"A7",X"03",X"06",
		X"FF",X"EE",X"DD",X"FF",X"EE",X"DD",X"CC",X"BB",X"AA",X"CC",X"BB",X"AA",X"99",X"88",X"77",X"99",
		X"88",X"77",X"00",X"00",X"30",X"07",X"00",X"2A",X"0C",X"01",X"72",X"2A",X"0A",X"01",X"00",X"30",
		X"07",X"07",X"81",X"30",X"05",X"07",X"00",X"54",X"30",X"02",X"00",X"60",X"0A",X"01",X"75",X"60",
		X"09",X"01",X"00",X"66",X"05",X"14",X"84",X"66",X"04",X"14",X"00",X"DE",X"30",X"05",X"02",X"05",
		X"08",X"00",X"08",X"00",X"88",X"80",X"08",X"00",X"80",X"80",X"02",X"05",X"55",X"50",X"50",X"50",
		X"55",X"50",X"05",X"00",X"05",X"00",X"02",X"05",X"66",X"60",X"60",X"60",X"66",X"60",X"06",X"00",
		X"06",X"00",X"64",X"03",X"2D",X"FA",X"A9",X"FF",X"01",X"FF",X"FA",X"2C",X"50",X"FA",X"AA",X"FF",
		X"01",X"FF",X"FA",X"28",X"2D",X"F0",X"B3",X"FF",X"01",X"FF",X"20",X"49",X"4E",X"46",X"45",X"52",
		X"4E",X"4F",X"20",X"28",X"43",X"29",X"20",X"31",X"39",X"38",X"34",X"20",X"57",X"49",X"4C",X"4C",
		X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",
		X"20",X"49",X"4E",X"43",X"2E",X"20",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"33",X"11",X"31",X"28",X"31",X"4C",X"64",X"EA",X"64",X"E1",X"7E",X"39",X"4D",X"7E",X"39",
		X"29",X"7E",X"39",X"2E",X"7E",X"39",X"33",X"7E",X"46",X"C4",X"7E",X"3B",X"45",X"7E",X"72",X"F6",
		X"7E",X"3C",X"52",X"7E",X"74",X"0C",X"7E",X"3C",X"65",X"00",X"00",X"00",X"00",X"12",X"15",X"00",
		X"00",X"00",X"01",X"25",X"20",X"00",X"21",X"20",X"34",X"40",X"00",X"A1",X"28",X"40",X"00",X"10",
		X"A0",X"23",X"53",X"31",X"10",X"A1",X"20",X"64",X"42",X"10",X"A1",X"20",X"74",X"40",X"01",X"A2",
		X"24",X"85",X"53",X"00",X"A2",X"28",X"A2",X"20",X"20",X"A0",X"23",X"9D",X"00",X"20",X"A2",X"25",
		X"24",X"42",X"20",X"A1",X"20",X"34",X"44",X"02",X"A2",X"24",X"45",X"53",X"00",X"A2",X"28",X"54",
		X"22",X"30",X"A0",X"23",X"60",X"D0",X"30",X"A2",X"26",X"71",X"A2",X"30",X"A1",X"20",X"84",X"44",
		X"02",X"A2",X"24",X"95",X"53",X"00",X"A2",X"28",X"A4",X"42",X"40",X"A0",X"23",X"90",X"0D",X"40",
		X"A2",X"27",X"64",X"44",X"40",X"A1",X"20",X"74",X"41",X"02",X"A2",X"24",X"85",X"53",X"00",X"A2",
		X"28",X"A4",X"40",X"40",X"A0",X"23",X"9D",X"00",X"40",X"A1",X"25",X"64",X"42",X"40",X"A1",X"20",
		X"74",X"46",X"02",X"A2",X"24",X"85",X"53",X"00",X"A2",X"28",X"A4",X"42",X"40",X"A0",X"23",X"90",
		X"D0",X"40",X"A1",X"26",X"64",X"44",X"40",X"AA",X"20",X"74",X"41",X"02",X"AA",X"24",X"85",X"53",
		X"00",X"AA",X"28",X"A4",X"40",X"40",X"A0",X"23",X"90",X"0D",X"40",X"A1",X"27",X"64",X"42",X"40",
		X"AA",X"20",X"74",X"46",X"02",X"AA",X"24",X"85",X"53",X"00",X"AA",X"28",X"A4",X"20",X"40",X"A0",
		X"23",X"9D",X"00",X"40",X"A1",X"25",X"64",X"44",X"40",X"AA",X"20",X"74",X"44",X"02",X"AA",X"24",
		X"85",X"53",X"00",X"AA",X"28",X"A4",X"40",X"40",X"A0",X"23",X"90",X"D0",X"40",X"A1",X"26",X"64",
		X"42",X"40",X"AA",X"20",X"74",X"46",X"02",X"AA",X"24",X"85",X"53",X"00",X"AA",X"28",X"A4",X"44",
		X"40",X"A0",X"23",X"F0",X"00",X"00",X"AA",X"00",X"68",X"B4",X"65",X"A5",X"00",X"04",X"01",X"3C",
		X"62",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"AC",X"05",X"20",X"90",X"2B",X"00",X"00",
		X"00",X"00",X"90",X"B7",X"01",X"FC",X"01",X"55",X"00",X"00",X"25",X"02",X"68",X"BD",X"65",X"B7",
		X"00",X"44",X"01",X"4C",X"62",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"BC",X"6C",X"20",
		X"90",X"3A",X"00",X"00",X"00",X"00",X"90",X"B8",X"02",X"FE",X"01",X"66",X"00",X"00",X"25",X"02",
		X"72",X"FD",X"6F",X"2F",X"00",X"84",X"01",X"5C",X"62",X"18",X"77",X"D8",X"77",X"CF",X"72",X"EE",
		X"6F",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"B7",X"03",X"FE",X"01",X"BB",
		X"10",X"02",X"05",X"02",X"73",X"74",X"70",X"26",X"00",X"C2",X"01",X"6C",X"62",X"18",X"77",X"DB",
		X"77",X"D2",X"73",X"65",X"6F",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"B8",
		X"03",X"FE",X"01",X"99",X"10",X"02",X"07",X"02",X"74",X"12",X"70",X"91",X"01",X"00",X"01",X"7C",
		X"62",X"18",X"77",X"DE",X"77",X"D5",X"74",X"0A",X"6F",X"16",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"B9",X"03",X"FE",X"01",X"FF",X"10",X"02",X"09",X"02",X"4E",X"4F",X"4D",X"99",
		X"02",X"46",X"02",X"5E",X"4B",X"64",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FE",X"03",X"00",X"08",X"02",X"12",X"02",
		X"45",X"F2",X"45",X"74",X"02",X"AE",X"02",X"CE",X"43",X"B7",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FE",X"01",X"00",
		X"00",X"00",X"20",X"02",X"60",X"56",X"60",X"56",X"03",X"02",X"03",X"12",X"61",X"D4",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"FE",X"01",X"00",X"00",X"00",X"15",X"02",X"77",X"F2",X"78",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"61",X"60",X"64",X"63",X"6F",X"70",X"71",X"A7",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"8E",X"5A",X"AD",X"86",X"01",X"5F",X"BD",X"E0",X"63",X"BD",
		X"33",X"0B",X"CC",X"31",X"28",X"ED",X"A8",X"22",X"86",X"04",X"34",X"02",X"7F",X"B8",X"35",X"34",
		X"20",X"1F",X"23",X"10",X"8E",X"66",X"E6",X"CC",X"01",X"00",X"BD",X"E0",X"78",X"BD",X"33",X"0B",
		X"35",X"10",X"10",X"AF",X"88",X"44",X"6F",X"A8",X"44",X"CC",X"31",X"28",X"ED",X"A8",X"22",X"B6",
		X"B8",X"35",X"26",X"04",X"10",X"BF",X"B8",X"35",X"6A",X"E4",X"26",X"D3",X"DE",X"21",X"35",X"82",
		X"10",X"8E",X"5A",X"AD",X"86",X"02",X"5F",X"BD",X"E0",X"63",X"BD",X"33",X"0B",X"CC",X"31",X"4C",
		X"ED",X"A8",X"22",X"86",X"04",X"34",X"02",X"7F",X"B8",X"37",X"34",X"20",X"1F",X"23",X"10",X"8E",
		X"66",X"E6",X"CC",X"02",X"00",X"BD",X"E0",X"78",X"BD",X"33",X"0B",X"35",X"10",X"10",X"AF",X"88",
		X"44",X"6F",X"A8",X"44",X"CC",X"31",X"4C",X"ED",X"A8",X"22",X"B6",X"B8",X"37",X"26",X"04",X"10",
		X"BF",X"B8",X"37",X"6A",X"E4",X"26",X"D3",X"DE",X"21",X"35",X"82",X"25",X"01",X"39",X"7E",X"E0",
		X"00",X"86",X"11",X"A7",X"51",X"A7",X"52",X"8E",X"31",X"23",X"96",X"68",X"2A",X"03",X"8E",X"30",
		X"2E",X"AF",X"48",X"0F",X"90",X"86",X"01",X"B7",X"DF",X"0F",X"CC",X"30",X"FF",X"BD",X"E0",X"66",
		X"96",X"90",X"34",X"02",X"BD",X"E0",X"AD",X"BD",X"11",X"20",X"4F",X"5F",X"DD",X"B7",X"97",X"B9",
		X"96",X"6D",X"26",X"16",X"10",X"8E",X"3A",X"0A",X"8E",X"10",X"F9",X"C6",X"11",X"A6",X"A0",X"27",
		X"09",X"88",X"7C",X"80",X"41",X"BD",X"E0",X"09",X"20",X"F3",X"A6",X"E0",X"2A",X"0C",X"EC",X"48",
		X"FD",X"B8",X"0C",X"CC",X"30",X"29",X"ED",X"48",X"20",X"10",X"86",X"01",X"9B",X"6D",X"19",X"97",
		X"6D",X"96",X"68",X"2A",X"05",X"C6",X"11",X"BD",X"3B",X"B1",X"C6",X"11",X"BD",X"3B",X"CC",X"AE",
		X"48",X"E6",X"04",X"54",X"54",X"54",X"C4",X"1E",X"27",X"09",X"8E",X"32",X"46",X"3A",X"AE",X"84",
		X"BD",X"E0",X"75",X"86",X"1E",X"B7",X"B7",X"78",X"8E",X"B7",X"79",X"10",X"8E",X"B8",X"3C",X"A6",
		X"A4",X"31",X"23",X"A7",X"80",X"8C",X"B7",X"82",X"23",X"F5",X"FC",X"B8",X"89",X"FD",X"B7",X"87",
		X"86",X"06",X"BD",X"E0",X"7D",X"AE",X"48",X"E6",X"84",X"54",X"54",X"54",X"54",X"A6",X"03",X"84",
		X"0F",X"BD",X"E0",X"99",X"18",X"00",X"05",X"86",X"01",X"BD",X"E0",X"7D",X"DC",X"6F",X"B3",X"E0",
		X"86",X"26",X"F4",X"7F",X"CB",X"60",X"10",X"8E",X"3F",X"88",X"86",X"30",X"C6",X"FF",X"BD",X"E0",
		X"63",X"FC",X"B8",X"14",X"26",X"0B",X"86",X"1E",X"BD",X"E0",X"7D",X"FC",X"D0",X"28",X"FD",X"D0",
		X"3E",X"CC",X"40",X"A7",X"DD",X"6F",X"86",X"01",X"97",X"28",X"86",X"04",X"97",X"71",X"97",X"72",
		X"CC",X"00",X"04",X"ED",X"C8",X"2F",X"FC",X"B8",X"14",X"27",X"1B",X"ED",X"C8",X"16",X"BD",X"69",
		X"26",X"EC",X"5A",X"44",X"56",X"1F",X"98",X"E6",X"5E",X"FD",X"B8",X"16",X"EC",X"4C",X"FD",X"B8",
		X"1D",X"EC",X"4E",X"FD",X"B8",X"1F",X"86",X"02",X"BD",X"E0",X"7D",X"5F",X"BD",X"3B",X"B1",X"BD",
		X"3B",X"CC",X"CC",X"01",X"FF",X"BD",X"E0",X"66",X"CC",X"02",X"FF",X"BD",X"E0",X"66",X"7C",X"B8",
		X"30",X"96",X"31",X"27",X"03",X"BD",X"32",X"75",X"96",X"40",X"27",X"03",X"BD",X"32",X"C0",X"86",
		X"02",X"BD",X"E0",X"7D",X"AE",X"48",X"A6",X"03",X"44",X"44",X"44",X"44",X"BD",X"39",X"4D",X"B6",
		X"B8",X"32",X"27",X"46",X"10",X"8E",X"38",X"99",X"86",X"0C",X"5F",X"BD",X"E0",X"63",X"34",X"01",
		X"1A",X"F0",X"7F",X"CB",X"A0",X"8E",X"03",X"24",X"86",X"05",X"BD",X"E0",X"83",X"1F",X"01",X"30",
		X"02",X"86",X"05",X"BD",X"E0",X"83",X"FD",X"C8",X"82",X"30",X"04",X"86",X"05",X"BD",X"E0",X"83",
		X"FD",X"C8",X"86",X"ED",X"28",X"F7",X"B8",X"31",X"CC",X"BE",X"1F",X"FD",X"C8",X"84",X"86",X"00",
		X"BD",X"E0",X"96",X"86",X"FF",X"B7",X"CB",X"A0",X"35",X"01",X"86",X"01",X"97",X"28",X"FC",X"B8",
		X"95",X"FD",X"B8",X"2A",X"FC",X"B8",X"98",X"FD",X"B8",X"2C",X"FC",X"B8",X"9B",X"FD",X"B8",X"2E",
		X"B6",X"B8",X"90",X"B7",X"B8",X"25",X"CC",X"01",X"C2",X"ED",X"C8",X"5C",X"FC",X"B8",X"0C",X"27",
		X"14",X"B6",X"B8",X"A2",X"F6",X"B8",X"A5",X"FD",X"B8",X"0E",X"B6",X"B8",X"A8",X"B7",X"B8",X"10",
		X"BD",X"38",X"77",X"20",X"47",X"B6",X"B8",X"32",X"27",X"03",X"BD",X"38",X"77",X"AE",X"48",X"A6",
		X"84",X"84",X"0F",X"B7",X"B8",X"0E",X"A6",X"01",X"44",X"44",X"44",X"44",X"B7",X"B8",X"0F",X"A6",
		X"01",X"84",X"0F",X"B7",X"B8",X"10",X"A6",X"02",X"44",X"44",X"44",X"44",X"B7",X"B8",X"11",X"A6",
		X"02",X"84",X"0F",X"B7",X"B8",X"12",X"96",X"31",X"27",X"53",X"96",X"40",X"27",X"4F",X"8E",X"B8",
		X"0E",X"86",X"4C",X"BD",X"3B",X"A0",X"BD",X"3B",X"A0",X"BD",X"3B",X"A0",X"B6",X"B8",X"10",X"BB",
		X"B8",X"0F",X"BB",X"B8",X"0E",X"80",X"0D",X"23",X"20",X"10",X"8E",X"B8",X"0E",X"8D",X"06",X"8D",
		X"04",X"8D",X"02",X"20",X"E7",X"E6",X"A0",X"27",X"0F",X"A1",X"3F",X"22",X"07",X"40",X"AB",X"3F",
		X"A7",X"3F",X"4F",X"39",X"A0",X"3F",X"6F",X"3F",X"39",X"8E",X"B8",X"11",X"86",X"80",X"BD",X"3B",
		X"A0",X"F6",X"B8",X"11",X"C1",X"04",X"23",X"05",X"C6",X"04",X"F7",X"B8",X"11",X"B6",X"B8",X"11",
		X"BB",X"B8",X"12",X"BB",X"B8",X"0E",X"BB",X"B8",X"0F",X"BB",X"B8",X"10",X"80",X"0D",X"23",X"0C",
		X"10",X"8E",X"B8",X"0E",X"8D",X"BF",X"8D",X"BD",X"8D",X"BB",X"20",X"E1",X"B6",X"B8",X"14",X"27",
		X"11",X"B6",X"B8",X"0E",X"BA",X"B8",X"0F",X"BA",X"B8",X"10",X"27",X"06",X"8E",X"78",X"0D",X"BD",
		X"E0",X"75",X"B6",X"B8",X"11",X"27",X"1A",X"10",X"8E",X"46",X"C4",X"86",X"04",X"C6",X"FF",X"BD",
		X"E0",X"63",X"BD",X"33",X"0B",X"0C",X"90",X"86",X"03",X"BD",X"E0",X"7D",X"7A",X"B8",X"11",X"26",
		X"E6",X"B6",X"B8",X"0E",X"27",X"0D",X"BD",X"39",X"29",X"86",X"03",X"BD",X"E0",X"7D",X"7A",X"B8",
		X"0E",X"26",X"F3",X"B6",X"B8",X"0F",X"27",X"0D",X"BD",X"39",X"2E",X"86",X"03",X"BD",X"E0",X"7D",
		X"7A",X"B8",X"0F",X"26",X"F3",X"B6",X"B8",X"10",X"27",X"0D",X"BD",X"39",X"33",X"86",X"03",X"BD",
		X"E0",X"7D",X"7A",X"B8",X"10",X"26",X"F3",X"10",X"8E",X"3B",X"FB",X"FC",X"B8",X"14",X"27",X"09",
		X"86",X"0F",X"B7",X"B8",X"23",X"10",X"8E",X"3C",X"65",X"CC",X"0F",X"FF",X"BD",X"E0",X"63",X"86",
		X"08",X"BD",X"E0",X"7D",X"B6",X"B8",X"12",X"27",X"0B",X"BD",X"3B",X"51",X"BD",X"33",X"0B",X"7A",
		X"B8",X"12",X"26",X"F5",X"B6",X"B8",X"66",X"B7",X"B7",X"82",X"96",X"68",X"10",X"2A",X"DB",X"08",
		X"BE",X"B8",X"0C",X"26",X"0C",X"AE",X"48",X"30",X"05",X"8C",X"31",X"23",X"25",X"03",X"8E",X"30",
		X"8D",X"AF",X"48",X"86",X"0B",X"A7",X"4A",X"A7",X"4B",X"6F",X"4C",X"86",X"01",X"BD",X"E0",X"7D",
		X"8E",X"B8",X"2A",X"EC",X"81",X"27",X"05",X"83",X"00",X"01",X"ED",X"1E",X"8C",X"B8",X"2E",X"23",
		X"F2",X"7A",X"B7",X"78",X"2E",X"2D",X"86",X"1E",X"B7",X"B7",X"78",X"8E",X"B7",X"7A",X"A6",X"80",
		X"27",X"02",X"6A",X"1F",X"8C",X"B7",X"7F",X"23",X"F5",X"B6",X"B8",X"34",X"26",X"15",X"FC",X"B7",
		X"7D",X"81",X"0A",X"25",X"02",X"86",X"0A",X"C1",X"0A",X"25",X"02",X"C6",X"0A",X"FD",X"B7",X"7D",
		X"7A",X"B8",X"34",X"B6",X"B8",X"14",X"27",X"26",X"B6",X"B8",X"22",X"27",X"24",X"B6",X"B8",X"21",
		X"27",X"1F",X"86",X"0B",X"A7",X"4A",X"A7",X"4B",X"6F",X"4C",X"CC",X"01",X"2C",X"7D",X"B8",X"24",
		X"27",X"03",X"CC",X"02",X"58",X"10",X"B3",X"B7",X"87",X"25",X"03",X"FD",X"B7",X"87",X"7E",X"37",
		X"2D",X"FC",X"B7",X"87",X"C3",X"FF",X"FF",X"2E",X"35",X"7C",X"B8",X"13",X"2A",X"03",X"7A",X"B8",
		X"13",X"B6",X"B8",X"84",X"B7",X"B7",X"80",X"B6",X"B8",X"87",X"B7",X"B7",X"81",X"86",X"FF",X"97",
		X"B5",X"BD",X"3B",X"45",X"25",X"1B",X"86",X"FF",X"B7",X"B8",X"22",X"FC",X"B8",X"89",X"C3",X"FF",
		X"EC",X"2E",X"03",X"FC",X"B8",X"89",X"10",X"83",X"00",X"5A",X"25",X"02",X"44",X"56",X"FD",X"B7",
		X"87",X"B6",X"B8",X"13",X"B1",X"B7",X"86",X"23",X"24",X"6A",X"4C",X"2E",X"20",X"86",X"1E",X"A7",
		X"4C",X"6A",X"4A",X"2E",X"18",X"BD",X"3B",X"45",X"25",X"0F",X"A6",X"4B",X"44",X"81",X"03",X"22",
		X"02",X"86",X"03",X"A7",X"4B",X"A7",X"4A",X"20",X"04",X"6F",X"4A",X"6F",X"4C",X"EC",X"C8",X"5C",
		X"C3",X"FF",X"FF",X"ED",X"C8",X"5C",X"26",X"0E",X"CC",X"01",X"2C",X"ED",X"C8",X"5C",X"7C",X"B8",
		X"25",X"2A",X"03",X"7A",X"B8",X"25",X"96",X"90",X"10",X"2E",X"FE",X"FF",X"7F",X"B8",X"30",X"BD",
		X"E0",X"A7",X"BD",X"39",X"FF",X"BD",X"3B",X"E7",X"CC",X"00",X"F0",X"BD",X"E0",X"66",X"0F",X"32",
		X"0F",X"41",X"86",X"02",X"BD",X"E0",X"7D",X"FC",X"B8",X"0C",X"26",X"06",X"96",X"90",X"10",X"27",
		X"00",X"F5",X"8E",X"77",X"F8",X"FC",X"B8",X"0C",X"27",X"03",X"8E",X"77",X"FE",X"BD",X"E0",X"75",
		X"86",X"02",X"BD",X"E0",X"7D",X"BD",X"E0",X"AA",X"BD",X"E0",X"AD",X"FC",X"B8",X"16",X"26",X"03",
		X"CC",X"48",X"2E",X"C3",X"FF",X"F8",X"FD",X"9A",X"4A",X"7C",X"DF",X"0F",X"B6",X"DF",X"0F",X"B7",
		X"9A",X"4E",X"0F",X"28",X"0C",X"2F",X"0C",X"3E",X"8E",X"11",X"1A",X"FC",X"B8",X"0C",X"27",X"12",
		X"7A",X"DF",X"0F",X"8E",X"11",X"44",X"7F",X"9A",X"4E",X"96",X"B7",X"91",X"B8",X"24",X"03",X"7C",
		X"9A",X"4E",X"AD",X"84",X"86",X"01",X"97",X"28",X"34",X"01",X"1A",X"F0",X"CC",X"1F",X"10",X"FD",
		X"C8",X"86",X"8E",X"05",X"10",X"BF",X"C8",X"84",X"CC",X"12",X"00",X"F7",X"C8",X"81",X"B7",X"C8",
		X"80",X"0D",X"49",X"27",X"09",X"8E",X"6C",X"10",X"BF",X"C8",X"84",X"B7",X"C8",X"80",X"35",X"01",
		X"FC",X"B8",X"0C",X"27",X"36",X"10",X"8E",X"31",X"28",X"BD",X"3A",X"36",X"0D",X"49",X"27",X"07",
		X"10",X"8E",X"31",X"4C",X"BD",X"3A",X"36",X"10",X"8E",X"31",X"28",X"BD",X"3A",X"E3",X"0D",X"49",
		X"27",X"07",X"10",X"8E",X"31",X"4C",X"BD",X"3A",X"E3",X"8E",X"78",X"01",X"BD",X"E0",X"75",X"FC",
		X"11",X"47",X"DD",X"6F",X"86",X"1B",X"BD",X"E0",X"7D",X"20",X"3C",X"86",X"05",X"BD",X"E0",X"7D",
		X"8E",X"77",X"FB",X"BD",X"E0",X"75",X"10",X"8E",X"31",X"28",X"96",X"90",X"43",X"27",X"04",X"10",
		X"8E",X"31",X"4C",X"10",X"AF",X"C8",X"22",X"86",X"1E",X"A7",X"C8",X"12",X"CC",X"01",X"02",X"BD",
		X"11",X"1D",X"8E",X"77",X"FE",X"12",X"12",X"12",X"86",X"01",X"BD",X"E0",X"7D",X"6A",X"C8",X"12",
		X"26",X"EA",X"86",X"03",X"BD",X"E0",X"7D",X"86",X"03",X"BD",X"E0",X"7D",X"BD",X"E0",X"AD",X"BD",
		X"11",X"23",X"0F",X"4C",X"7E",X"33",X"2A",X"4F",X"5F",X"FD",X"B8",X"2A",X"FD",X"B8",X"2C",X"FD",
		X"B8",X"2E",X"FD",X"B7",X"7D",X"F7",X"B7",X"7F",X"86",X"99",X"B7",X"B8",X"25",X"86",X"01",X"B7",
		X"B7",X"83",X"B7",X"B7",X"84",X"B7",X"B7",X"85",X"39",X"6F",X"4A",X"B6",X"B8",X"9F",X"A7",X"4B",
		X"86",X"01",X"BD",X"E0",X"7D",X"A6",X"4A",X"E6",X"48",X"3D",X"C3",X"BE",X"1F",X"1F",X"01",X"C6",
		X"07",X"10",X"8E",X"39",X"1B",X"6A",X"4B",X"27",X"2C",X"A6",X"A0",X"30",X"86",X"A6",X"84",X"85",
		X"F0",X"27",X"08",X"8B",X"10",X"85",X"F0",X"26",X"02",X"8B",X"10",X"A7",X"84",X"A6",X"A0",X"30",
		X"86",X"A6",X"84",X"85",X"0F",X"27",X"07",X"4C",X"85",X"0F",X"26",X"02",X"8B",X"F1",X"A7",X"80",
		X"5A",X"26",X"D6",X"20",X"BB",X"B6",X"B8",X"33",X"27",X"B1",X"34",X"10",X"8E",X"77",X"C3",X"BD",
		X"E0",X"9E",X"35",X"10",X"A6",X"A0",X"30",X"86",X"A6",X"84",X"84",X"0F",X"A7",X"84",X"A6",X"A0",
		X"30",X"86",X"A6",X"84",X"84",X"F0",X"A7",X"80",X"5A",X"26",X"E9",X"6C",X"4A",X"7A",X"B8",X"31",
		X"26",X"89",X"8E",X"77",X"C6",X"BD",X"E0",X"9E",X"7E",X"E0",X"69",X"E4",X"07",X"07",X"07",X"00",
		X"07",X"00",X"00",X"F9",X"00",X"F9",X"F9",X"F9",X"00",X"8E",X"31",X"70",X"20",X"08",X"8E",X"31",
		X"94",X"20",X"03",X"8E",X"31",X"B8",X"10",X"8E",X"55",X"C0",X"86",X"03",X"C6",X"FF",X"BD",X"E0",
		X"63",X"BD",X"33",X"0B",X"AF",X"A8",X"22",X"0C",X"90",X"7C",X"B8",X"34",X"39",X"34",X"02",X"10",
		X"8E",X"39",X"F5",X"8E",X"B7",X"89",X"E6",X"A0",X"E7",X"05",X"E7",X"0B",X"30",X"0C",X"8C",X"B7",
		X"FB",X"25",X"F3",X"CC",X"00",X"04",X"ED",X"C8",X"2F",X"A6",X"E4",X"27",X"63",X"34",X"02",X"10",
		X"8E",X"B7",X"89",X"8E",X"00",X"41",X"A6",X"89",X"9A",X"42",X"26",X"4B",X"A6",X"89",X"90",X"C1",
		X"26",X"45",X"A6",X"89",X"91",X"02",X"2F",X"3F",X"84",X"0F",X"81",X"01",X"27",X"0C",X"81",X"02",
		X"27",X"08",X"81",X"04",X"27",X"04",X"81",X"08",X"26",X"2D",X"BD",X"5F",X"B1",X"27",X"28",X"34",
		X"10",X"1F",X"10",X"F3",X"91",X"00",X"58",X"49",X"58",X"49",X"54",X"54",X"ED",X"C8",X"16",X"8D",
		X"21",X"EC",X"C8",X"16",X"1E",X"89",X"ED",X"C8",X"16",X"8D",X"17",X"35",X"10",X"6A",X"E4",X"2F",
		X"0D",X"10",X"8C",X"B7",X"FB",X"22",X"07",X"30",X"01",X"8C",X"09",X"40",X"25",X"A8",X"35",X"02",
		X"35",X"82",X"BD",X"69",X"26",X"AE",X"C8",X"14",X"86",X"81",X"A7",X"89",X"90",X"C1",X"AF",X"A4",
		X"EC",X"5A",X"44",X"56",X"86",X"1A",X"24",X"02",X"8A",X"20",X"A7",X"24",X"1F",X"98",X"E6",X"5E",
		X"ED",X"22",X"31",X"26",X"39",X"22",X"55",X"66",X"77",X"99",X"BB",X"EE",X"44",X"AA",X"DD",X"8E",
		X"B7",X"89",X"6F",X"80",X"8C",X"B8",X"01",X"25",X"F9",X"39",X"37",X"28",X"25",X"2D",X"2C",X"21",
		X"25",X"26",X"37",X"17",X"32",X"10",X"37",X"3E",X"36",X"35",X"39",X"37",X"1E",X"28",X"2B",X"2B",
		X"28",X"30",X"24",X"22",X"37",X"2C",X"2B",X"2C",X"32",X"23",X"21",X"26",X"25",X"28",X"32",X"22",
		X"37",X"28",X"25",X"32",X"13",X"00",X"AE",X"A8",X"12",X"86",X"00",X"BD",X"E0",X"83",X"10",X"83",
		X"77",X"77",X"10",X"27",X"00",X"9C",X"34",X"01",X"1A",X"F0",X"BF",X"C8",X"84",X"CC",X"1F",X"30",
		X"FD",X"C8",X"86",X"CC",X"12",X"77",X"F7",X"C8",X"81",X"B7",X"C8",X"80",X"86",X"03",X"B7",X"BF",
		X"FF",X"B7",X"C8",X"00",X"4F",X"5F",X"FD",X"80",X"EE",X"86",X"01",X"B7",X"BF",X"FF",X"B7",X"C8",
		X"00",X"35",X"01",X"E6",X"A8",X"1F",X"34",X"16",X"A6",X"B8",X"1A",X"1C",X"DE",X"19",X"A7",X"E4",
		X"AE",X"62",X"30",X"89",X"06",X"04",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"BD",X"E0",X"2C",X"CC",
		X"A8",X"44",X"BD",X"E0",X"25",X"CC",X"A9",X"44",X"AE",X"62",X"30",X"89",X"05",X"0C",X"BD",X"E0",
		X"25",X"CC",X"AA",X"44",X"AE",X"62",X"30",X"89",X"02",X"14",X"BD",X"E0",X"25",X"AE",X"62",X"30",
		X"89",X"06",X"1C",X"EC",X"E4",X"AB",X"E4",X"19",X"AB",X"E4",X"19",X"85",X"F0",X"26",X"02",X"8A",
		X"F0",X"BD",X"E0",X"17",X"86",X"2D",X"BD",X"E0",X"09",X"86",X"00",X"BD",X"E0",X"09",X"BD",X"E0",
		X"09",X"BD",X"E0",X"09",X"AE",X"62",X"30",X"89",X"02",X"26",X"CC",X"6E",X"44",X"BD",X"E0",X"25",
		X"35",X"16",X"39",X"BD",X"3A",X"36",X"A6",X"B8",X"1A",X"C6",X"03",X"DE",X"21",X"10",X"AF",X"C8",
		X"22",X"20",X"00",X"ED",X"C8",X"3E",X"EC",X"E1",X"ED",X"C8",X"44",X"86",X"04",X"BD",X"E0",X"7D",
		X"EC",X"C8",X"3E",X"85",X"0F",X"27",X"10",X"6A",X"C8",X"3E",X"86",X"03",X"BD",X"11",X"1D",X"8E",
		X"77",X"54",X"BD",X"E0",X"75",X"20",X"E4",X"5C",X"6E",X"D8",X"44",X"ED",X"C8",X"3E",X"EC",X"E1",
		X"ED",X"C8",X"44",X"86",X"04",X"BD",X"E0",X"7D",X"EC",X"C8",X"3E",X"85",X"F0",X"27",X"12",X"80",
		X"10",X"A7",X"C8",X"3E",X"86",X"03",X"BD",X"11",X"1D",X"8E",X"77",X"54",X"BD",X"E0",X"75",X"20",
		X"E2",X"5C",X"6E",X"D8",X"44",X"8D",X"0A",X"25",X"07",X"86",X"FF",X"A7",X"A8",X"4B",X"1C",X"FE",
		X"39",X"B6",X"B8",X"23",X"43",X"85",X"0C",X"27",X"44",X"F6",X"B7",X"86",X"C1",X"03",X"24",X"3D",
		X"10",X"8E",X"41",X"12",X"86",X"05",X"5F",X"BD",X"E0",X"63",X"25",X"31",X"6F",X"A8",X"4B",X"7C",
		X"B7",X"86",X"CC",X"32",X"00",X"ED",X"A8",X"22",X"F6",X"B8",X"23",X"C4",X"0C",X"27",X"04",X"C8",
		X"0C",X"20",X"0E",X"C6",X"04",X"86",X"80",X"B8",X"B8",X"23",X"B7",X"B8",X"23",X"2B",X"02",X"C6",
		X"08",X"E7",X"A8",X"4E",X"FA",X"B8",X"23",X"F7",X"B8",X"23",X"1C",X"FE",X"39",X"1A",X"01",X"39",
		X"34",X"02",X"E6",X"84",X"27",X"09",X"3D",X"4D",X"26",X"01",X"4C",X"AB",X"84",X"A7",X"80",X"35",
		X"82",X"86",X"62",X"8E",X"3D",X"70",X"BD",X"E0",X"10",X"30",X"89",X"03",X"00",X"96",X"6D",X"85",
		X"F0",X"26",X"06",X"30",X"89",X"FD",X"00",X"8A",X"F0",X"7E",X"E0",X"17",X"AE",X"48",X"A6",X"04",
		X"84",X"0F",X"27",X"12",X"8E",X"32",X"65",X"A6",X"86",X"81",X"A7",X"26",X"03",X"7C",X"B8",X"32",
		X"8E",X"00",X"80",X"7E",X"E0",X"56",X"39",X"96",X"31",X"9A",X"40",X"27",X"01",X"39",X"10",X"8E",
		X"11",X"2C",X"86",X"31",X"5F",X"BD",X"E0",X"63",X"7E",X"E0",X"69",X"8E",X"77",X"F5",X"BD",X"E0",
		X"9E",X"BD",X"E0",X"99",X"EF",X"DA",X"05",X"BD",X"E0",X"99",X"EF",X"DD",X"05",X"25",X"08",X"8E",
		X"3C",X"07",X"86",X"01",X"7E",X"E0",X"6C",X"8E",X"90",X"02",X"AE",X"84",X"2A",X"F1",X"A6",X"11",
		X"81",X"03",X"26",X"F6",X"A6",X"88",X"51",X"27",X"F1",X"34",X"10",X"6F",X"88",X"51",X"10",X"AE",
		X"88",X"22",X"CC",X"76",X"C9",X"ED",X"88",X"25",X"EC",X"A8",X"10",X"ED",X"88",X"27",X"FC",X"EF",
		X"CA",X"ED",X"88",X"58",X"86",X"0C",X"A7",X"88",X"5C",X"AE",X"2A",X"BD",X"E0",X"75",X"35",X"10",
		X"20",X"C8",X"34",X"10",X"BE",X"B8",X"18",X"A7",X"84",X"E7",X"88",X"10",X"EC",X"E4",X"A7",X"01",
		X"E7",X"88",X"11",X"35",X"90",X"86",X"05",X"A7",X"48",X"CC",X"7F",X"7F",X"FD",X"B7",X"3E",X"7F",
		X"B7",X"43",X"7F",X"B7",X"47",X"86",X"04",X"BD",X"E0",X"7D",X"CC",X"1B",X"9B",X"8E",X"1C",X"9C",
		X"BD",X"3C",X"52",X"86",X"01",X"BD",X"E0",X"7D",X"CC",X"19",X"99",X"8E",X"1A",X"9A",X"BD",X"3C",
		X"52",X"BD",X"3F",X"7C",X"10",X"23",X"00",X"9E",X"86",X"02",X"BD",X"E0",X"7D",X"86",X"F0",X"B4",
		X"B8",X"23",X"B7",X"B8",X"23",X"BD",X"3F",X"26",X"25",X"55",X"2F",X"27",X"BD",X"3F",X"16",X"CC",
		X"22",X"23",X"BD",X"3D",X"9C",X"26",X"6E",X"86",X"04",X"BD",X"E0",X"7D",X"CC",X"22",X"23",X"BD",
		X"3D",X"9C",X"26",X"61",X"BD",X"3F",X"7C",X"23",X"6D",X"BD",X"3F",X"3B",X"BD",X"3F",X"26",X"25",
		X"2E",X"2E",X"E9",X"BD",X"3F",X"16",X"CC",X"A3",X"A2",X"BD",X"3D",X"9C",X"26",X"47",X"86",X"04",
		X"BD",X"E0",X"7D",X"CC",X"A3",X"A2",X"BD",X"3D",X"9C",X"26",X"3A",X"BD",X"3F",X"7C",X"23",X"46",
		X"BD",X"3F",X"3B",X"BD",X"3F",X"26",X"25",X"07",X"2F",X"E9",X"20",X"B0",X"BD",X"3F",X"16",X"CC",
		X"19",X"99",X"BD",X"3D",X"9C",X"26",X"1E",X"86",X"04",X"BD",X"E0",X"7D",X"CC",X"19",X"99",X"BD",
		X"3D",X"9C",X"26",X"11",X"BD",X"3F",X"7C",X"23",X"1D",X"BD",X"3F",X"3B",X"BD",X"3F",X"26",X"25",
		X"EB",X"2E",X"8C",X"20",X"B1",X"BD",X"3F",X"16",X"86",X"04",X"BD",X"E0",X"7D",X"B6",X"B8",X"23",
		X"84",X"0C",X"26",X"F4",X"20",X"C9",X"86",X"0F",X"BA",X"B8",X"23",X"B7",X"B8",X"23",X"CC",X"19",
		X"99",X"8E",X"1A",X"9A",X"BD",X"3C",X"52",X"86",X"01",X"BD",X"E0",X"7D",X"CC",X"1B",X"9B",X"8E",
		X"1C",X"9C",X"BD",X"3C",X"52",X"86",X"02",X"BD",X"E0",X"7D",X"CC",X"1D",X"9D",X"8E",X"1E",X"9E",
		X"BD",X"3C",X"52",X"86",X"01",X"BD",X"E0",X"7D",X"8E",X"3F",X"10",X"AF",X"4D",X"AF",X"4F",X"EC",
		X"84",X"10",X"BE",X"B8",X"18",X"E7",X"C8",X"11",X"E7",X"C8",X"12",X"A7",X"21",X"88",X"80",X"A7",
		X"A8",X"11",X"ED",X"C8",X"13",X"4F",X"A7",X"C8",X"15",X"A7",X"C8",X"16",X"BD",X"3D",X"B6",X"86",
		X"06",X"BD",X"E0",X"7D",X"EC",X"C8",X"13",X"26",X"F3",X"7E",X"3C",X"75",X"7D",X"B8",X"21",X"27",
		X"08",X"CC",X"1B",X"9B",X"8E",X"1C",X"9C",X"20",X"03",X"8E",X"1A",X"9A",X"BD",X"3C",X"52",X"B6",
		X"B8",X"23",X"84",X"0C",X"39",X"09",X"10",X"BE",X"B8",X"18",X"AE",X"4D",X"B6",X"B7",X"3E",X"B1",
		X"3D",X"B5",X"22",X"2D",X"8C",X"3F",X"14",X"26",X"09",X"8E",X"77",X"E7",X"BD",X"E0",X"75",X"7E",
		X"3E",X"60",X"A6",X"C8",X"15",X"26",X"0D",X"6A",X"C8",X"15",X"34",X"10",X"8E",X"77",X"E4",X"BD",
		X"E0",X"75",X"35",X"10",X"6A",X"C8",X"11",X"2E",X"77",X"30",X"02",X"EC",X"84",X"8D",X"44",X"20",
		X"6F",X"6F",X"C8",X"13",X"8C",X"3F",X"10",X"27",X"67",X"A6",X"C8",X"15",X"27",X"0D",X"6F",X"C8",
		X"15",X"34",X"10",X"8E",X"77",X"EA",X"BD",X"E0",X"75",X"35",X"10",X"6C",X"C8",X"13",X"6A",X"C8",
		X"11",X"2E",X"4D",X"7F",X"B7",X"43",X"BE",X"B8",X"1B",X"86",X"F6",X"A4",X"89",X"91",X"03",X"A7",
		X"89",X"91",X"03",X"A7",X"89",X"91",X"04",X"A7",X"89",X"91",X"05",X"AE",X"4D",X"EC",X"83",X"8D",
		X"02",X"20",X"2D",X"A7",X"21",X"E7",X"C8",X"11",X"E7",X"C8",X"13",X"AF",X"4D",X"8C",X"3F",X"14",
		X"26",X"1D",X"86",X"03",X"A7",X"C8",X"11",X"B7",X"B7",X"43",X"BE",X"B8",X"1B",X"86",X"09",X"AA",
		X"89",X"91",X"03",X"A7",X"89",X"91",X"03",X"A7",X"89",X"91",X"04",X"A7",X"89",X"91",X"05",X"39",
		X"AE",X"4F",X"B6",X"B7",X"3F",X"B1",X"3D",X"B5",X"22",X"2D",X"8C",X"3F",X"14",X"26",X"09",X"8E",
		X"77",X"E7",X"BD",X"E0",X"75",X"7E",X"3F",X"09",X"A6",X"C8",X"16",X"26",X"0D",X"6A",X"C8",X"16",
		X"34",X"10",X"8E",X"77",X"E4",X"BD",X"E0",X"75",X"35",X"10",X"6A",X"C8",X"12",X"2E",X"7A",X"30",
		X"02",X"EC",X"84",X"8D",X"44",X"20",X"72",X"6F",X"C8",X"14",X"8C",X"3F",X"10",X"27",X"6A",X"A6",
		X"C8",X"16",X"27",X"0D",X"6F",X"C8",X"16",X"34",X"10",X"8E",X"77",X"EA",X"BD",X"E0",X"75",X"35",
		X"10",X"6C",X"C8",X"14",X"6A",X"C8",X"12",X"2E",X"50",X"7F",X"B7",X"47",X"BE",X"B8",X"1B",X"86",
		X"F9",X"A4",X"89",X"91",X"42",X"A7",X"89",X"91",X"42",X"A7",X"89",X"91",X"82",X"A7",X"89",X"91",
		X"C2",X"AE",X"4F",X"EC",X"83",X"8D",X"02",X"20",X"30",X"88",X"80",X"A7",X"A8",X"11",X"E7",X"C8",
		X"12",X"E7",X"C8",X"14",X"AF",X"4F",X"8C",X"3F",X"14",X"26",X"1D",X"86",X"03",X"A7",X"C8",X"12",
		X"B7",X"B7",X"47",X"BE",X"B8",X"1B",X"86",X"06",X"AA",X"89",X"91",X"42",X"A7",X"89",X"91",X"42",
		X"A7",X"89",X"91",X"82",X"A7",X"89",X"91",X"C2",X"39",X"CC",X"7F",X"7F",X"FD",X"B7",X"3E",X"39",
		X"1E",X"01",X"1F",X"01",X"20",X"0A",X"CC",X"19",X"99",X"BE",X"B8",X"18",X"A7",X"84",X"E7",X"88",
		X"10",X"86",X"04",X"7E",X"E0",X"7D",X"FC",X"B7",X"3C",X"26",X"03",X"1A",X"01",X"39",X"34",X"02",
		X"7F",X"B7",X"3C",X"7F",X"B7",X"3D",X"E1",X"E0",X"1C",X"FE",X"39",X"6A",X"48",X"26",X"38",X"BD",
		X"E0",X"72",X"49",X"C6",X"1E",X"3D",X"8B",X"07",X"24",X"02",X"86",X"FF",X"A7",X"48",X"BE",X"B8",
		X"18",X"A6",X"84",X"E6",X"88",X"10",X"ED",X"4B",X"EC",X"E1",X"ED",X"49",X"CC",X"21",X"A1",X"A7",
		X"84",X"E7",X"88",X"10",X"86",X"02",X"BD",X"E0",X"7D",X"EC",X"4B",X"BE",X"B8",X"18",X"A7",X"84",
		X"E7",X"88",X"10",X"EC",X"49",X"34",X"06",X"86",X"04",X"7E",X"E0",X"7D",X"FC",X"B7",X"3E",X"B1",
		X"3D",X"B5",X"23",X"03",X"F1",X"3D",X"B5",X"39",X"CC",X"40",X"53",X"ED",X"48",X"86",X"01",X"A7",
		X"4A",X"A7",X"4B",X"8E",X"40",X"53",X"AF",X"48",X"8E",X"40",X"86",X"AF",X"4C",X"6F",X"4E",X"6F",
		X"4F",X"6F",X"C8",X"10",X"8D",X"32",X"B6",X"B8",X"14",X"27",X"25",X"8D",X"43",X"B6",X"B8",X"AA",
		X"27",X"1E",X"96",X"6D",X"81",X"30",X"25",X"18",X"BD",X"E0",X"72",X"34",X"02",X"C6",X"2F",X"3D",
		X"1F",X"01",X"35",X"02",X"C6",X"60",X"3D",X"30",X"86",X"86",X"90",X"5F",X"30",X"8B",X"6C",X"84",
		X"8E",X"3F",X"A4",X"86",X"01",X"7E",X"E0",X"6C",X"6A",X"4A",X"2E",X"13",X"AE",X"48",X"EC",X"81",
		X"FD",X"D0",X"50",X"A6",X"80",X"2A",X"04",X"40",X"8E",X"40",X"53",X"AF",X"48",X"A7",X"4A",X"39",
		X"6A",X"4B",X"2E",X"17",X"86",X"07",X"97",X"72",X"AE",X"4C",X"EC",X"81",X"FD",X"D0",X"5E",X"A6",
		X"80",X"2A",X"04",X"40",X"8E",X"40",X"86",X"AF",X"4C",X"A7",X"4B",X"FC",X"D0",X"5E",X"FD",X"D0",
		X"5C",X"FD",X"D0",X"56",X"FD",X"D0",X"46",X"6A",X"4E",X"2E",X"0F",X"BD",X"E0",X"72",X"84",X"0F",
		X"8B",X"0A",X"A7",X"4E",X"CC",X"FF",X"FF",X"FD",X"D0",X"56",X"6A",X"4F",X"2A",X"0F",X"BD",X"E0",
		X"72",X"84",X"07",X"8B",X"0A",X"A7",X"4F",X"CC",X"FF",X"FF",X"FD",X"D0",X"46",X"6A",X"C8",X"10",
		X"2A",X"10",X"BD",X"E0",X"72",X"84",X"07",X"8B",X"0A",X"A7",X"C8",X"10",X"CC",X"FF",X"FF",X"FD",
		X"D0",X"5C",X"39",X"0F",X"D0",X"02",X"0F",X"B0",X"02",X"0F",X"A0",X"02",X"0F",X"80",X"02",X"0F",
		X"60",X"02",X"0F",X"80",X"02",X"0F",X"A0",X"02",X"0F",X"80",X"02",X"0F",X"60",X"02",X"0F",X"40",
		X"02",X"00",X"00",X"04",X"F0",X"4F",X"04",X"F0",X"8F",X"04",X"F0",X"BF",X"04",X"F0",X"8F",X"04",
		X"F0",X"4F",X"04",X"00",X"00",X"FC",X"0F",X"D0",X"06",X"0F",X"B0",X"02",X"0F",X"A0",X"02",X"0F",
		X"80",X"02",X"0F",X"60",X"04",X"0F",X"80",X"02",X"0F",X"A0",X"02",X"0F",X"80",X"02",X"0F",X"70",
		X"02",X"0F",X"50",X"02",X"0F",X"30",X"FC",X"FC",X"D0",X"5E",X"FD",X"81",X"3E",X"FC",X"D0",X"56",
		X"FD",X"81",X"36",X"FC",X"D0",X"5C",X"FD",X"81",X"3C",X"FC",X"D0",X"46",X"FD",X"81",X"26",X"B6",
		X"B8",X"14",X"26",X"1B",X"FC",X"D0",X"3E",X"FD",X"81",X"1E",X"FD",X"81",X"3E",X"FD",X"81",X"5E",
		X"FD",X"81",X"7E",X"FD",X"81",X"9E",X"FD",X"81",X"BE",X"FD",X"81",X"DE",X"FD",X"81",X"FE",X"0A",
		X"71",X"2A",X"2E",X"86",X"04",X"97",X"71",X"FC",X"81",X"50",X"FD",X"81",X"30",X"FC",X"81",X"70",
		X"FD",X"81",X"50",X"FC",X"81",X"90",X"FD",X"81",X"70",X"FC",X"81",X"B0",X"FD",X"81",X"90",X"FC",
		X"81",X"D0",X"FD",X"81",X"B0",X"FC",X"81",X"F0",X"FD",X"81",X"D0",X"FC",X"D0",X"50",X"FD",X"81",
		X"F0",X"39",X"6F",X"C8",X"5E",X"C6",X"04",X"E7",X"C8",X"20",X"B6",X"B8",X"1A",X"A7",X"42",X"BE",
		X"B8",X"14",X"26",X"03",X"8E",X"10",X"10",X"10",X"8E",X"42",X"9D",X"A6",X"C8",X"4E",X"85",X"04",
		X"26",X"04",X"10",X"8E",X"42",X"A5",X"EC",X"A1",X"30",X"8B",X"AF",X"C8",X"16",X"CC",X"0C",X"0C",
		X"ED",X"C8",X"54",X"86",X"08",X"A7",X"C8",X"56",X"CC",X"01",X"01",X"ED",X"4A",X"6F",X"C8",X"11",
		X"34",X"20",X"BD",X"54",X"1F",X"35",X"20",X"B6",X"B8",X"66",X"A7",X"C8",X"3B",X"EC",X"5A",X"E3",
		X"A4",X"ED",X"5A",X"E6",X"42",X"E7",X"C8",X"46",X"CB",X"17",X"E7",X"42",X"EC",X"5D",X"83",X"00",
		X"17",X"E3",X"22",X"ED",X"5D",X"A6",X"23",X"E6",X"21",X"40",X"50",X"ED",X"C8",X"4F",X"6F",X"43",
		X"6F",X"C8",X"12",X"FC",X"EF",X"C2",X"ED",X"C8",X"5A",X"AE",X"24",X"AF",X"C8",X"29",X"CC",X"02",
		X"05",X"ED",X"C8",X"1E",X"BE",X"B8",X"18",X"27",X"40",X"8E",X"77",X"7E",X"BD",X"6A",X"33",X"86",
		X"0A",X"BD",X"E0",X"7D",X"BD",X"42",X"54",X"BE",X"B8",X"18",X"86",X"21",X"E6",X"C8",X"4E",X"C5",
		X"08",X"26",X"05",X"88",X"80",X"30",X"88",X"10",X"A7",X"84",X"A6",X"5E",X"A7",X"5F",X"6F",X"5E",
		X"86",X"03",X"BD",X"E0",X"7D",X"BD",X"42",X"54",X"A6",X"5F",X"A7",X"5E",X"6A",X"C8",X"1E",X"2E",
		X"CE",X"86",X"14",X"BD",X"E0",X"7D",X"BD",X"42",X"54",X"8E",X"77",X"84",X"BD",X"6A",X"33",X"AE",
		X"C8",X"29",X"30",X"02",X"AF",X"C8",X"29",X"8D",X"74",X"86",X"08",X"BD",X"E0",X"7D",X"8D",X"64",
		X"8D",X"6B",X"25",X"09",X"86",X"01",X"BD",X"E0",X"7D",X"8D",X"59",X"20",X"F3",X"86",X"04",X"BD",
		X"E0",X"7D",X"86",X"04",X"BD",X"E0",X"7D",X"8D",X"4B",X"AE",X"C8",X"29",X"30",X"02",X"AF",X"C8",
		X"29",X"6A",X"C8",X"1F",X"26",X"EC",X"FC",X"EF",X"BC",X"ED",X"C8",X"5A",X"4F",X"5F",X"ED",X"C8",
		X"47",X"ED",X"C8",X"37",X"86",X"01",X"A7",X"C8",X"45",X"EC",X"C8",X"16",X"ED",X"C8",X"1C",X"ED",
		X"C8",X"1A",X"CC",X"04",X"04",X"ED",X"C8",X"1E",X"A6",X"C8",X"4E",X"43",X"B4",X"B8",X"23",X"B7",
		X"B8",X"23",X"C6",X"08",X"BD",X"45",X"36",X"8D",X"0B",X"6A",X"C8",X"1F",X"26",X"F4",X"BD",X"45",
		X"35",X"7E",X"42",X"AD",X"B6",X"B8",X"21",X"27",X"03",X"A7",X"C8",X"5E",X"39",X"EC",X"C8",X"4F",
		X"27",X"38",X"81",X"02",X"23",X"02",X"86",X"02",X"34",X"02",X"40",X"AB",X"C8",X"4F",X"A7",X"C8",
		X"4F",X"35",X"02",X"AB",X"5E",X"A7",X"5E",X"1D",X"2B",X"08",X"C1",X"03",X"2F",X"0A",X"C6",X"03",
		X"20",X"06",X"C1",X"FD",X"2C",X"02",X"C6",X"FD",X"34",X"04",X"50",X"EB",X"C8",X"50",X"E7",X"C8",
		X"50",X"35",X"04",X"E3",X"5A",X"ED",X"5A",X"1C",X"FE",X"39",X"1A",X"01",X"39",X"09",X"00",X"FF",
		X"D5",X"FF",X"F1",X"02",X"DE",X"00",X"09",X"00",X"2A",X"FF",X"F1",X"02",X"EA",X"86",X"07",X"A7",
		X"C8",X"39",X"EC",X"C8",X"16",X"BD",X"44",X"7B",X"4F",X"5F",X"ED",X"C8",X"33",X"A7",X"5F",X"A7",
		X"C8",X"18",X"86",X"0F",X"A7",X"C8",X"24",X"8E",X"77",X"78",X"BD",X"44",X"41",X"AD",X"D8",X"25",
		X"AD",X"D8",X"27",X"E6",X"43",X"10",X"27",X"00",X"D0",X"E7",X"C8",X"20",X"8E",X"64",X"E1",X"E6",
		X"85",X"8E",X"64",X"EA",X"3A",X"1F",X"12",X"EC",X"24",X"E3",X"C8",X"14",X"1F",X"01",X"EC",X"26",
		X"E3",X"C8",X"16",X"BD",X"44",X"CA",X"24",X"10",X"A6",X"43",X"43",X"A4",X"C8",X"24",X"26",X"02",
		X"86",X"0F",X"A7",X"C8",X"24",X"7E",X"43",X"A9",X"34",X"06",X"BD",X"45",X"0F",X"35",X"06",X"BD",
		X"44",X"7B",X"86",X"0F",X"A7",X"C8",X"24",X"10",X"8E",X"77",X"90",X"BD",X"44",X"16",X"27",X"61",
		X"25",X"04",X"10",X"8E",X"77",X"8A",X"1F",X"21",X"BD",X"44",X"41",X"BD",X"45",X"26",X"BD",X"68",
		X"49",X"25",X"45",X"A6",X"C8",X"4B",X"26",X"08",X"BD",X"45",X"26",X"BD",X"68",X"49",X"25",X"38",
		X"BD",X"44",X"16",X"26",X"E6",X"A6",X"C8",X"4B",X"26",X"31",X"C6",X"08",X"E7",X"C8",X"4D",X"E6",
		X"5F",X"57",X"E7",X"5F",X"27",X"25",X"E6",X"C8",X"4D",X"BD",X"45",X"36",X"BD",X"68",X"49",X"25",
		X"17",X"BD",X"44",X"4A",X"26",X"F0",X"6F",X"C8",X"4D",X"BD",X"45",X"35",X"BD",X"68",X"49",X"25",
		X"07",X"BD",X"44",X"16",X"26",X"F3",X"20",X"D7",X"7E",X"43",X"B7",X"8E",X"77",X"78",X"BD",X"44",
		X"41",X"6A",X"C8",X"13",X"E6",X"43",X"BD",X"72",X"8D",X"BD",X"45",X"35",X"BD",X"68",X"49",X"25",
		X"26",X"BD",X"45",X"45",X"BD",X"68",X"49",X"25",X"1E",X"E6",X"43",X"BD",X"72",X"B6",X"6F",X"C8",
		X"13",X"BD",X"45",X"45",X"BD",X"68",X"49",X"25",X"0E",X"6F",X"C8",X"13",X"BD",X"45",X"45",X"BD",
		X"68",X"49",X"25",X"03",X"7E",X"42",X"CD",X"1F",X"12",X"7A",X"B7",X"86",X"2E",X"06",X"8E",X"77",
		X"96",X"BD",X"E0",X"9E",X"CC",X"01",X"01",X"ED",X"C8",X"18",X"A6",X"A8",X"10",X"A7",X"C8",X"10",
		X"FC",X"EF",X"D8",X"ED",X"C8",X"5A",X"BD",X"44",X"61",X"AE",X"C8",X"22",X"1E",X"23",X"EC",X"88",
		X"22",X"BD",X"11",X"1D",X"8E",X"77",X"A5",X"BD",X"E0",X"75",X"DE",X"21",X"BD",X"45",X"45",X"A6",
		X"C8",X"18",X"2E",X"F8",X"6F",X"5E",X"86",X"01",X"BD",X"E0",X"7D",X"7E",X"E0",X"69",X"BD",X"44",
		X"61",X"6F",X"5E",X"7A",X"B7",X"86",X"2E",X"06",X"8E",X"77",X"96",X"BD",X"E0",X"9E",X"86",X"01",
		X"BD",X"E0",X"7D",X"7E",X"E0",X"69",X"A6",X"C8",X"46",X"8B",X"17",X"A1",X"42",X"34",X"01",X"27",
		X"1E",X"25",X"0E",X"8E",X"77",X"8A",X"BD",X"44",X"41",X"6C",X"42",X"6A",X"5E",X"6A",X"5F",X"20",
		X"0C",X"8E",X"77",X"90",X"BD",X"44",X"41",X"6A",X"42",X"6C",X"5E",X"6C",X"5F",X"A6",X"5F",X"35",
		X"81",X"96",X"B5",X"27",X"02",X"30",X"03",X"7E",X"E0",X"9E",X"A6",X"5F",X"27",X"12",X"2A",X"08",
		X"6C",X"42",X"6A",X"5E",X"6C",X"5F",X"20",X"06",X"6A",X"42",X"6C",X"5E",X"6A",X"5F",X"1C",X"FE",
		X"39",X"34",X"10",X"8E",X"B8",X"04",X"EC",X"C8",X"31",X"10",X"A3",X"84",X"26",X"04",X"6F",X"84",
		X"6F",X"01",X"30",X"02",X"8C",X"B8",X"0A",X"23",X"F0",X"35",X"90",X"AE",X"C8",X"16",X"ED",X"C8",
		X"31",X"BC",X"B8",X"04",X"26",X"04",X"FD",X"B8",X"04",X"39",X"BC",X"B8",X"06",X"26",X"04",X"FD",
		X"B8",X"06",X"39",X"BC",X"B8",X"08",X"26",X"04",X"FD",X"B8",X"08",X"39",X"BC",X"B8",X"0A",X"26",
		X"04",X"FD",X"B8",X"0A",X"39",X"BE",X"B8",X"04",X"26",X"04",X"FD",X"B8",X"04",X"39",X"BE",X"B8",
		X"06",X"26",X"04",X"FD",X"B8",X"06",X"39",X"BE",X"B8",X"08",X"26",X"04",X"FD",X"B8",X"08",X"39",
		X"BE",X"B8",X"0A",X"26",X"04",X"FD",X"B8",X"0A",X"39",X"39",X"34",X"10",X"8E",X"B8",X"04",X"8D",
		X"14",X"25",X"10",X"27",X"0E",X"8D",X"0E",X"25",X"0A",X"27",X"08",X"8D",X"08",X"25",X"04",X"27",
		X"02",X"8D",X"02",X"35",X"90",X"34",X"06",X"6D",X"84",X"27",X"1E",X"A0",X"84",X"24",X"01",X"40",
		X"81",X"02",X"24",X"15",X"E0",X"01",X"24",X"01",X"50",X"C1",X"02",X"24",X"0C",X"EC",X"C8",X"16",
		X"10",X"A3",X"84",X"27",X"06",X"1A",X"01",X"35",X"86",X"30",X"02",X"1C",X"FE",X"35",X"86",X"8C",
		X"09",X"40",X"24",X"11",X"A6",X"89",X"91",X"02",X"2B",X"0B",X"85",X"0F",X"27",X"07",X"44",X"44",
		X"84",X"38",X"A7",X"C8",X"46",X"39",X"C6",X"08",X"A6",X"5F",X"2A",X"01",X"40",X"81",X"04",X"25",
		X"02",X"C6",X"10",X"20",X"01",X"5F",X"A6",X"C8",X"20",X"8E",X"64",X"BD",X"EB",X"86",X"AE",X"C8",
		X"2F",X"3A",X"AF",X"C8",X"29",X"A6",X"C8",X"12",X"27",X"03",X"6A",X"C8",X"12",X"E6",X"C8",X"1E",
		X"C0",X"02",X"2A",X"02",X"C6",X"04",X"E7",X"C8",X"1E",X"AE",X"C8",X"2D",X"3A",X"AF",X"C8",X"2B",
		X"BD",X"E0",X"88",X"86",X"01",X"7E",X"E0",X"7D",X"EC",X"C8",X"16",X"ED",X"C8",X"47",X"86",X"1E",
		X"A7",X"C8",X"12",X"39",X"AE",X"D8",X"37",X"2A",X"EF",X"EC",X"C8",X"33",X"27",X"EA",X"A6",X"88",
		X"51",X"27",X"E5",X"AE",X"C8",X"14",X"8C",X"09",X"40",X"24",X"E8",X"A6",X"89",X"91",X"02",X"2F",
		X"E2",X"BD",X"5F",X"B1",X"27",X"DD",X"AE",X"D8",X"37",X"EC",X"88",X"16",X"A0",X"C8",X"16",X"2A",
		X"01",X"40",X"E0",X"C8",X"17",X"2A",X"01",X"50",X"34",X"02",X"E1",X"E4",X"25",X"02",X"E7",X"E4",
		X"35",X"02",X"B1",X"B7",X"80",X"22",X"3A",X"EC",X"C8",X"16",X"A3",X"C8",X"47",X"27",X"17",X"4D",
		X"2A",X"01",X"40",X"5D",X"2A",X"01",X"50",X"34",X"04",X"A1",X"E4",X"22",X"02",X"A6",X"E4",X"35",
		X"04",X"B1",X"B7",X"81",X"22",X"05",X"A6",X"C8",X"12",X"2E",X"16",X"BD",X"69",X"A2",X"25",X"11",
		X"54",X"E7",X"C8",X"12",X"54",X"EB",X"C8",X"12",X"E7",X"C8",X"12",X"EC",X"C8",X"16",X"ED",X"C8",
		X"47",X"39",X"A6",X"C8",X"4B",X"27",X"0A",X"B6",X"B8",X"21",X"26",X"64",X"A6",X"C8",X"5E",X"26",
		X"5F",X"B6",X"B7",X"73",X"26",X"0B",X"A6",X"C8",X"3B",X"BD",X"6E",X"53",X"EC",X"C8",X"33",X"26",
		X"03",X"6F",X"43",X"39",X"6A",X"C8",X"45",X"2E",X"38",X"BD",X"75",X"32",X"A7",X"C8",X"45",X"44",
		X"44",X"AB",X"C8",X"45",X"A7",X"C8",X"45",X"26",X"07",X"86",X"0A",X"A7",X"C8",X"45",X"20",X"E1",
		X"E6",X"80",X"E5",X"C8",X"24",X"26",X"17",X"E6",X"80",X"E5",X"C8",X"24",X"26",X"10",X"E6",X"80",
		X"E5",X"C8",X"24",X"26",X"09",X"E6",X"80",X"E5",X"C8",X"24",X"26",X"02",X"20",X"C3",X"E7",X"43",
		X"39",X"EC",X"5A",X"2B",X"C4",X"10",X"83",X"01",X"20",X"24",X"BE",X"A6",X"5D",X"26",X"BA",X"39",
		X"CC",X"46",X"6C",X"ED",X"C8",X"25",X"CC",X"46",X"8D",X"ED",X"C8",X"27",X"A6",X"C8",X"20",X"85",
		X"0C",X"26",X"02",X"48",X"48",X"A7",X"43",X"EC",X"5A",X"10",X"83",X"01",X"20",X"22",X"0B",X"A6",
		X"5E",X"81",X"20",X"22",X"04",X"81",X"10",X"22",X"01",X"39",X"7E",X"43",X"FE",X"A6",X"43",X"27",
		X"03",X"A7",X"C8",X"21",X"39",X"34",X"16",X"A6",X"C8",X"3A",X"27",X"11",X"6F",X"C8",X"3A",X"7A",
		X"B8",X"02",X"2E",X"09",X"7F",X"B8",X"02",X"8E",X"77",X"AB",X"BD",X"E0",X"9E",X"35",X"96",X"34",
		X"16",X"A6",X"C8",X"3A",X"26",X"0C",X"6C",X"C8",X"3A",X"7C",X"B8",X"02",X"8E",X"77",X"A8",X"BD",
		X"E0",X"9E",X"35",X"96",X"7C",X"B8",X"24",X"8E",X"90",X"95",X"A6",X"81",X"2B",X"FC",X"EF",X"83",
		X"CC",X"31",X"DC",X"ED",X"C8",X"22",X"96",X"68",X"2B",X"0A",X"CC",X"95",X"58",X"B3",X"91",X"00",
		X"1F",X"01",X"20",X"05",X"BD",X"54",X"90",X"30",X"1E",X"30",X"02",X"EC",X"81",X"26",X"08",X"9C",
		X"62",X"25",X"F8",X"9E",X"60",X"20",X"F4",X"4D",X"26",X"04",X"1F",X"98",X"30",X"01",X"30",X"1E",
		X"4D",X"2B",X"E6",X"85",X"F0",X"27",X"E2",X"85",X"10",X"26",X"DE",X"85",X"0F",X"27",X"DA",X"A6",
		X"89",X"09",X"40",X"26",X"D4",X"CC",X"02",X"52",X"ED",X"C8",X"29",X"C6",X"02",X"A6",X"88",X"40",
		X"2F",X"41",X"85",X"10",X"26",X"3D",X"A6",X"89",X"09",X"80",X"26",X"37",X"A6",X"88",X"C0",X"2F",
		X"32",X"85",X"10",X"26",X"2E",X"A6",X"89",X"09",X"00",X"26",X"28",X"E7",X"C8",X"20",X"BD",X"55",
		X"68",X"AE",X"C8",X"14",X"30",X"88",X"C0",X"AF",X"C8",X"4B",X"30",X"89",X"00",X"80",X"AF",X"C8",
		X"4D",X"CC",X"18",X"0C",X"ED",X"C8",X"54",X"86",X"08",X"A7",X"C8",X"56",X"CC",X"01",X"00",X"ED",
		X"4A",X"20",X"4E",X"CC",X"02",X"48",X"ED",X"C8",X"29",X"C6",X"01",X"A6",X"01",X"10",X"2F",X"FF",
		X"78",X"85",X"10",X"10",X"26",X"FF",X"72",X"A6",X"89",X"09",X"41",X"10",X"26",X"FF",X"6A",X"A6",
		X"1F",X"10",X"2F",X"FF",X"64",X"85",X"10",X"10",X"26",X"FF",X"5E",X"A6",X"89",X"09",X"3F",X"10",
		X"26",X"FF",X"56",X"E7",X"C8",X"20",X"BD",X"55",X"68",X"AE",X"C8",X"14",X"30",X"1F",X"AF",X"C8",
		X"4B",X"30",X"02",X"AF",X"C8",X"4D",X"CC",X"0C",X"18",X"ED",X"C8",X"54",X"CC",X"00",X"01",X"ED",
		X"4A",X"BD",X"53",X"FD",X"6F",X"C8",X"3A",X"BD",X"46",X"95",X"FC",X"EF",X"D2",X"ED",X"C8",X"5A",
		X"86",X"FF",X"A7",X"C8",X"5E",X"A6",X"C8",X"20",X"A7",X"C8",X"21",X"6F",X"C8",X"1E",X"6F",X"43",
		X"6F",X"C8",X"3F",X"6F",X"C8",X"40",X"6F",X"C8",X"43",X"6F",X"C8",X"3E",X"6F",X"C8",X"12",X"BD",
		X"4A",X"EB",X"EC",X"C8",X"16",X"E3",X"4A",X"ED",X"C8",X"1C",X"EC",X"C8",X"16",X"A3",X"4A",X"ED",
		X"C8",X"1A",X"6F",X"C8",X"18",X"C6",X"02",X"E7",X"C8",X"57",X"A6",X"43",X"27",X"06",X"A7",X"C8",
		X"20",X"BD",X"4A",X"EB",X"AD",X"D8",X"27",X"AD",X"D8",X"25",X"A6",X"43",X"27",X"1E",X"BD",X"49",
		X"D6",X"A6",X"89",X"9A",X"42",X"27",X"40",X"85",X"F0",X"27",X"25",X"A6",X"43",X"43",X"A4",X"C8",
		X"24",X"BD",X"49",X"AE",X"A7",X"C8",X"24",X"26",X"03",X"BD",X"4A",X"EB",X"7E",X"48",X"9F",X"A6",
		X"43",X"BD",X"49",X"AE",X"6A",X"C8",X"3B",X"2E",X"66",X"C6",X"03",X"E7",X"C8",X"3B",X"20",X"DD",
		X"81",X"02",X"22",X"EB",X"27",X"07",X"7D",X"B7",X"16",X"2A",X"D0",X"20",X"05",X"7D",X"B7",X"18",
		X"2A",X"C9",X"B6",X"B7",X"73",X"26",X"C4",X"86",X"0A",X"A7",X"C8",X"3B",X"AF",X"C8",X"31",X"BD",
		X"46",X"AF",X"BD",X"4A",X"1F",X"26",X"44",X"A6",X"C8",X"11",X"AA",X"89",X"9A",X"42",X"A7",X"89",
		X"9A",X"42",X"6A",X"C8",X"13",X"E6",X"43",X"BD",X"72",X"8D",X"AE",X"C8",X"31",X"BD",X"49",X"C1",
		X"BD",X"4A",X"80",X"BD",X"4A",X"40",X"AE",X"C8",X"31",X"BD",X"49",X"C1",X"AD",X"D8",X"27",X"6F",
		X"C8",X"13",X"BD",X"4A",X"80",X"A6",X"43",X"27",X"03",X"A7",X"C8",X"3F",X"7E",X"47",X"FA",X"6F",
		X"C8",X"13",X"BD",X"46",X"95",X"BD",X"4A",X"80",X"7E",X"47",X"FA",X"8E",X"77",X"3F",X"A6",X"43",
		X"E6",X"86",X"53",X"8E",X"64",X"E1",X"E6",X"85",X"8E",X"64",X"EA",X"3A",X"EC",X"04",X"E3",X"C8",
		X"14",X"1F",X"01",X"A6",X"89",X"9A",X"42",X"27",X"1D",X"85",X"F0",X"27",X"15",X"A6",X"43",X"43",
		X"A4",X"C8",X"24",X"A7",X"C8",X"24",X"10",X"26",X"FF",X"2D",X"BD",X"4A",X"EB",X"BD",X"49",X"AE",
		X"20",X"BD",X"81",X"02",X"22",X"F7",X"A6",X"C8",X"11",X"AA",X"89",X"9A",X"42",X"A7",X"89",X"9A",
		X"42",X"AF",X"C8",X"4F",X"AE",X"C8",X"31",X"A6",X"C8",X"11",X"AA",X"89",X"9A",X"42",X"A7",X"89",
		X"9A",X"42",X"BD",X"4A",X"7E",X"AD",X"D8",X"27",X"A6",X"43",X"AA",X"C8",X"20",X"8E",X"4A",X"0F",
		X"E6",X"86",X"BD",X"4A",X"AD",X"AD",X"D8",X"27",X"A6",X"43",X"A7",X"C8",X"20",X"BD",X"4A",X"7E",
		X"AD",X"D8",X"27",X"EC",X"C8",X"54",X"1E",X"89",X"ED",X"C8",X"54",X"EC",X"4A",X"1E",X"89",X"ED",
		X"4A",X"EC",X"C8",X"16",X"E3",X"4A",X"ED",X"C8",X"1C",X"EC",X"C8",X"16",X"A3",X"4A",X"ED",X"C8",
		X"1A",X"AE",X"C8",X"4B",X"A6",X"C8",X"11",X"43",X"A4",X"89",X"9A",X"42",X"A7",X"89",X"9A",X"42",
		X"AE",X"C8",X"31",X"AF",X"C8",X"4B",X"BD",X"49",X"C1",X"AE",X"C8",X"4D",X"A6",X"C8",X"11",X"43",
		X"A4",X"89",X"9A",X"42",X"A7",X"89",X"9A",X"42",X"AE",X"C8",X"4F",X"AF",X"C8",X"4D",X"BD",X"49",
		X"C1",X"A6",X"43",X"A7",X"C8",X"20",X"BD",X"4A",X"80",X"AD",X"D8",X"27",X"BD",X"4A",X"7E",X"7E",
		X"47",X"FA",X"20",X"49",X"4E",X"46",X"45",X"52",X"4E",X"4F",X"20",X"28",X"43",X"29",X"20",X"31",
		X"39",X"38",X"34",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",X"34",X"16",
		X"A6",X"43",X"27",X"0B",X"8E",X"77",X"3F",X"E6",X"86",X"53",X"E7",X"C8",X"3F",X"6F",X"43",X"35",
		X"96",X"E6",X"89",X"9A",X"42",X"C4",X"0F",X"27",X"0C",X"C1",X"02",X"22",X"08",X"B6",X"B7",X"73",
		X"26",X"03",X"7E",X"51",X"84",X"39",X"AE",X"C8",X"14",X"E6",X"C8",X"20",X"C5",X"09",X"27",X"17",
		X"81",X"04",X"23",X"03",X"30",X"02",X"39",X"26",X"04",X"30",X"88",X"40",X"39",X"44",X"25",X"04",
		X"30",X"88",X"C0",X"39",X"30",X"1E",X"39",X"81",X"04",X"23",X"03",X"30",X"01",X"39",X"26",X"05",
		X"30",X"89",X"00",X"80",X"39",X"44",X"25",X"04",X"30",X"88",X"80",X"39",X"30",X"1F",X"39",X"00",
		X"00",X"00",X"16",X"00",X"14",X"00",X"00",X"00",X"00",X"14",X"00",X"16",X"00",X"00",X"00",X"A6",
		X"C8",X"20",X"A1",X"43",X"27",X"19",X"10",X"8E",X"77",X"3F",X"E6",X"A6",X"E4",X"43",X"26",X"0F",
		X"EC",X"C8",X"4D",X"10",X"AE",X"C8",X"4B",X"10",X"AF",X"C8",X"4D",X"ED",X"C8",X"4B",X"4F",X"39",
		X"AE",X"C8",X"4D",X"27",X"0C",X"A6",X"C8",X"11",X"43",X"A4",X"89",X"9A",X"42",X"A7",X"89",X"9A",
		X"42",X"EC",X"C8",X"14",X"ED",X"C8",X"4D",X"EC",X"C8",X"4B",X"ED",X"C8",X"14",X"EC",X"C8",X"31",
		X"ED",X"C8",X"4B",X"E6",X"43",X"BD",X"72",X"8D",X"EC",X"06",X"E3",X"C8",X"16",X"ED",X"C8",X"16",
		X"E3",X"4A",X"ED",X"C8",X"1C",X"EC",X"C8",X"16",X"A3",X"4A",X"ED",X"C8",X"1A",X"39",X"20",X"3B",
		X"5F",X"A6",X"C8",X"51",X"85",X"02",X"27",X"33",X"E6",X"C8",X"1E",X"A6",X"43",X"27",X"2C",X"CB",
		X"02",X"85",X"03",X"26",X"08",X"C0",X"04",X"2A",X"09",X"C6",X"06",X"20",X"05",X"C1",X"06",X"23",
		X"01",X"5F",X"E7",X"C8",X"1E",X"CB",X"02",X"85",X"09",X"26",X"02",X"CB",X"0A",X"A6",X"C8",X"51",
		X"85",X"02",X"27",X"07",X"8E",X"02",X"46",X"3A",X"AF",X"C8",X"29",X"A6",X"C8",X"51",X"85",X"01",
		X"27",X"0F",X"8E",X"64",X"C6",X"A6",X"C8",X"21",X"E6",X"86",X"8E",X"02",X"5E",X"3A",X"AF",X"C8",
		X"2B",X"A6",X"C8",X"57",X"26",X"05",X"BD",X"E0",X"88",X"20",X"03",X"BD",X"E0",X"8B",X"86",X"01",
		X"E6",X"C8",X"51",X"C5",X"01",X"27",X"01",X"4C",X"7E",X"E0",X"7D",X"AE",X"C8",X"14",X"E6",X"89",
		X"91",X"02",X"BC",X"B7",X"49",X"27",X"1B",X"BC",X"B7",X"50",X"27",X"1B",X"BC",X"B7",X"57",X"27",
		X"1B",X"BC",X"B7",X"5E",X"27",X"1B",X"BC",X"B7",X"65",X"27",X"1B",X"BC",X"B7",X"6C",X"27",X"1B",
		X"20",X"1C",X"F6",X"B7",X"4B",X"20",X"17",X"F6",X"B7",X"52",X"20",X"12",X"F6",X"B7",X"59",X"20",
		X"0D",X"F6",X"B7",X"60",X"20",X"08",X"F6",X"B7",X"67",X"20",X"03",X"F6",X"B7",X"6E",X"C4",X"0F",
		X"A6",X"89",X"91",X"03",X"2F",X"06",X"85",X"10",X"27",X"02",X"C4",X"F7",X"A6",X"89",X"91",X"42",
		X"2F",X"06",X"85",X"10",X"27",X"02",X"C4",X"FB",X"A6",X"89",X"90",X"C2",X"2F",X"06",X"85",X"10",
		X"27",X"02",X"C4",X"FD",X"A6",X"89",X"91",X"01",X"2F",X"06",X"85",X"10",X"27",X"02",X"C4",X"FE",
		X"E7",X"C8",X"24",X"39",X"3F",X"20",X"FD",X"BD",X"46",X"95",X"CC",X"4B",X"AC",X"ED",X"C8",X"25",
		X"AE",X"C8",X"4B",X"A6",X"C8",X"11",X"43",X"1F",X"89",X"A4",X"89",X"9A",X"42",X"A7",X"89",X"9A",
		X"42",X"AE",X"C8",X"4D",X"E4",X"89",X"9A",X"42",X"E7",X"89",X"9A",X"42",X"CC",X"0C",X"0C",X"ED",
		X"C8",X"54",X"4F",X"5F",X"ED",X"4A",X"EC",X"C8",X"16",X"ED",X"C8",X"1C",X"ED",X"C8",X"1A",X"EB",
		X"C8",X"14",X"E7",X"48",X"6F",X"C8",X"57",X"6F",X"49",X"BD",X"4B",X"E3",X"A6",X"C8",X"51",X"27",
		X"03",X"6F",X"43",X"39",X"A6",X"C8",X"18",X"26",X"F8",X"6F",X"5E",X"AE",X"C8",X"14",X"A6",X"C8",
		X"11",X"43",X"A4",X"89",X"9A",X"42",X"A7",X"89",X"9A",X"42",X"0A",X"90",X"E6",X"C8",X"11",X"BD",
		X"51",X"50",X"CC",X"00",X"00",X"ED",X"84",X"BD",X"4B",X"E3",X"BD",X"46",X"95",X"7A",X"B8",X"24",
		X"7E",X"E0",X"69",X"8E",X"90",X"93",X"30",X"02",X"8C",X"90",X"9B",X"22",X"10",X"11",X"A3",X"84",
		X"26",X"F4",X"EC",X"02",X"ED",X"81",X"8C",X"90",X"9B",X"25",X"F7",X"6F",X"83",X"39",X"39",X"86",
		X"01",X"A7",X"C8",X"42",X"86",X"A0",X"A7",X"C8",X"41",X"CC",X"4C",X"0F",X"ED",X"C8",X"25",X"6A",
		X"C8",X"42",X"26",X"34",X"6F",X"43",X"CC",X"4C",X"28",X"ED",X"C8",X"25",X"BD",X"E0",X"72",X"C6",
		X"0F",X"3D",X"8B",X"0A",X"A7",X"C8",X"42",X"39",X"6F",X"43",X"6A",X"C8",X"41",X"26",X"03",X"6C",
		X"C8",X"41",X"6A",X"C8",X"42",X"26",X"F0",X"BD",X"E0",X"72",X"C6",X"3C",X"3D",X"8B",X"1E",X"A7",
		X"C8",X"42",X"CC",X"4C",X"0F",X"ED",X"C8",X"25",X"A6",X"C8",X"3F",X"8E",X"77",X"3F",X"A6",X"86",
		X"6A",X"C8",X"41",X"26",X"12",X"34",X"02",X"BD",X"E0",X"72",X"C6",X"1E",X"3D",X"8B",X"3C",X"A7",
		X"C8",X"42",X"35",X"02",X"43",X"20",X"14",X"A4",X"C8",X"24",X"26",X"08",X"A6",X"C8",X"3F",X"A6",
		X"86",X"43",X"20",X"07",X"8E",X"77",X"2F",X"E6",X"86",X"2A",X"03",X"A7",X"43",X"39",X"34",X"02",
		X"8E",X"4C",X"9B",X"E6",X"86",X"BD",X"E0",X"72",X"49",X"3D",X"1F",X"89",X"86",X"10",X"44",X"A5",
		X"E4",X"27",X"FB",X"E0",X"86",X"22",X"F7",X"35",X"04",X"20",X"E0",X"00",X"1E",X"3C",X"5A",X"1E",
		X"3C",X"5A",X"78",X"3C",X"5A",X"78",X"96",X"5A",X"78",X"96",X"B4",X"EC",X"A8",X"16",X"A0",X"C8",
		X"16",X"2A",X"01",X"40",X"E0",X"C8",X"17",X"2A",X"01",X"50",X"34",X"02",X"E1",X"E4",X"25",X"02",
		X"E7",X"E4",X"EC",X"88",X"16",X"A0",X"C8",X"16",X"2A",X"01",X"40",X"E0",X"C8",X"17",X"2A",X"01",
		X"50",X"34",X"02",X"E1",X"E0",X"22",X"02",X"1F",X"89",X"E1",X"E0",X"25",X"02",X"1E",X"12",X"39",
		X"F6",X"B7",X"73",X"27",X"06",X"96",X"68",X"10",X"2B",X"00",X"88",X"6A",X"C8",X"39",X"2E",X"1F",
		X"A7",X"C8",X"39",X"10",X"BE",X"B7",X"16",X"27",X"05",X"A6",X"A8",X"51",X"26",X"1C",X"BE",X"B7",
		X"18",X"27",X"05",X"A6",X"88",X"51",X"26",X"33",X"4F",X"5F",X"ED",X"C8",X"33",X"20",X"63",X"AE",
		X"D8",X"37",X"2A",X"F4",X"A6",X"88",X"51",X"27",X"EF",X"39",X"BE",X"B7",X"18",X"27",X"1A",X"A6",
		X"88",X"51",X"27",X"15",X"86",X"08",X"AB",X"42",X"A0",X"22",X"2B",X"0F",X"C6",X"08",X"EB",X"42",
		X"E0",X"02",X"2B",X"11",X"BD",X"4C",X"AB",X"20",X"0E",X"1E",X"12",X"86",X"08",X"AB",X"42",X"A0",
		X"02",X"2B",X"C5",X"20",X"02",X"1E",X"12",X"A6",X"02",X"A7",X"C8",X"35",X"A6",X"88",X"3A",X"A7",
		X"C8",X"36",X"EC",X"88",X"16",X"10",X"A3",X"C8",X"33",X"27",X"03",X"6C",X"C8",X"40",X"ED",X"C8",
		X"33",X"10",X"8E",X"B7",X"18",X"BC",X"B7",X"18",X"27",X"04",X"10",X"8E",X"B7",X"16",X"10",X"AF",
		X"C8",X"37",X"39",X"6F",X"C8",X"39",X"CC",X"6F",X"14",X"ED",X"C8",X"37",X"BE",X"B7",X"74",X"2A",
		X"87",X"CC",X"B7",X"74",X"ED",X"C8",X"37",X"A6",X"02",X"A7",X"C8",X"35",X"A6",X"88",X"3A",X"A7",
		X"C8",X"36",X"EC",X"88",X"16",X"ED",X"C8",X"33",X"39",X"B6",X"B8",X"63",X"BD",X"4C",X"E0",X"EC",
		X"C8",X"33",X"26",X"22",X"86",X"1E",X"A7",X"C8",X"12",X"A6",X"43",X"27",X"05",X"A1",X"C8",X"21",
		X"26",X"06",X"C6",X"05",X"E7",X"C8",X"43",X"39",X"6A",X"C8",X"43",X"2E",X"08",X"8D",X"F3",X"A7",
		X"C8",X"21",X"A7",X"C8",X"10",X"39",X"A6",X"C8",X"12",X"2F",X"03",X"6A",X"C8",X"12",X"A6",X"C8",
		X"3E",X"2F",X"03",X"6A",X"C8",X"3E",X"A6",X"C8",X"12",X"26",X"21",X"BD",X"71",X"72",X"25",X"C4",
		X"8D",X"37",X"27",X"09",X"E7",X"C8",X"12",X"27",X"04",X"81",X"0C",X"23",X"0F",X"81",X"3C",X"22",
		X"0C",X"BD",X"6A",X"C3",X"25",X"06",X"F6",X"B8",X"7B",X"E7",X"C8",X"12",X"39",X"A6",X"C8",X"12",
		X"2E",X"FA",X"A6",X"C8",X"3E",X"2E",X"F5",X"BD",X"6A",X"C3",X"25",X"F0",X"F6",X"B8",X"7E",X"E7",
		X"C8",X"3E",X"F6",X"B8",X"7B",X"E7",X"C8",X"12",X"39",X"34",X"02",X"E6",X"C8",X"21",X"A6",X"C8",
		X"10",X"E7",X"C8",X"10",X"F6",X"B8",X"8D",X"A1",X"C8",X"21",X"35",X"82",X"EC",X"C8",X"33",X"8E",
		X"76",X"CF",X"A0",X"C8",X"16",X"2A",X"04",X"40",X"30",X"88",X"10",X"E0",X"C8",X"17",X"2A",X"03",
		X"50",X"30",X"08",X"34",X"02",X"E1",X"E0",X"23",X"03",X"30",X"04",X"39",X"1E",X"89",X"39",X"A6",
		X"C8",X"24",X"27",X"27",X"E6",X"C8",X"40",X"27",X"15",X"E6",X"C8",X"3F",X"8E",X"77",X"3F",X"A4",
		X"85",X"26",X"0E",X"E6",X"C8",X"3F",X"8E",X"77",X"3F",X"A6",X"85",X"43",X"20",X"0D",X"A7",X"C8",
		X"40",X"8E",X"77",X"2F",X"E6",X"86",X"2B",X"03",X"BD",X"4E",X"7E",X"A7",X"43",X"39",X"85",X"0F",
		X"27",X"59",X"34",X"02",X"EC",X"C8",X"33",X"8E",X"76",X"CF",X"A0",X"C8",X"16",X"2A",X"04",X"40",
		X"30",X"88",X"10",X"E0",X"C8",X"17",X"2A",X"03",X"50",X"30",X"08",X"34",X"02",X"E1",X"E4",X"25",
		X"18",X"E7",X"E4",X"30",X"04",X"C1",X"0A",X"25",X"22",X"48",X"34",X"04",X"A1",X"E0",X"23",X"1B",
		X"BD",X"E0",X"72",X"24",X"16",X"30",X"1C",X"20",X"12",X"81",X"0A",X"25",X"0E",X"58",X"34",X"04",
		X"A1",X"E0",X"24",X"07",X"BD",X"E0",X"72",X"24",X"02",X"30",X"04",X"35",X"06",X"E5",X"80",X"26",
		X"14",X"E5",X"80",X"26",X"10",X"E5",X"80",X"26",X"03",X"A6",X"84",X"39",X"E5",X"84",X"27",X"05",
		X"BD",X"E0",X"72",X"25",X"F4",X"A6",X"82",X"39",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"13",X"21",X"17",X"E1",X"02",X"0B",X"04",X"0B",X"00",X"FF",X"04",X"12",X"20",X"16",X"C1",X"02",
		X"37",X"0A",X"63",X"02",X"08",X"01",X"01",X"01",X"35",X"81",X"06",X"37",X"0C",X"8F",X"04",X"09",
		X"01",X"01",X"01",X"32",X"C1",X"02",X"37",X"0A",X"63",X"04",X"FC",X"01",X"0F",X"1D",X"13",X"E1",
		X"06",X"0B",X"08",X"0B",X"00",X"FB",X"FC",X"0A",X"18",X"12",X"C1",X"06",X"37",X"0C",X"63",X"02",
		X"04",X"01",X"01",X"01",X"31",X"81",X"02",X"37",X"0A",X"8F",X"04",X"05",X"01",X"01",X"01",X"2E",
		X"C1",X"06",X"37",X"0C",X"63",X"04",X"F8",X"F9",X"07",X"15",X"0F",X"11",X"02",X"00",X"02",X"00",
		X"00",X"F7",X"F8",X"06",X"14",X"0E",X"01",X"00",X"00",X"00",X"00",X"02",X"00",X"FD",X"FD",X"FD",
		X"01",X"11",X"22",X"00",X"22",X"00",X"02",X"2B",X"FC",X"FC",X"FC",X"23",X"01",X"00",X"00",X"00",
		X"00",X"04",X"00",X"F8",X"F8",X"F8",X"01",X"11",X"22",X"00",X"22",X"00",X"04",X"27",X"F7",X"F7",
		X"F7",X"24",X"02",X"0E",X"00",X"0E",X"00",X"00",X"00",X"F3",X"01",X"25",X"1D",X"E2",X"10",X"16",
		X"12",X"16",X"00",X"FF",X"F6",X"04",X"24",X"20",X"C2",X"10",X"42",X"18",X"6E",X"0A",X"08",X"01",
		X"01",X"19",X"01",X"82",X"14",X"42",X"1A",X"9A",X"0C",X"09",X"01",X"01",X"16",X"01",X"C2",X"10",
		X"42",X"18",X"6E",X"0C",X"FC",X"F3",X"01",X"21",X"1D",X"E2",X"14",X"16",X"16",X"16",X"00",X"FB",
		X"EE",X"FC",X"20",X"18",X"C2",X"14",X"42",X"1A",X"6E",X"0A",X"04",X"05",X"01",X"15",X"01",X"82",
		X"10",X"42",X"18",X"9A",X"0C",X"05",X"01",X"01",X"12",X"01",X"C2",X"14",X"42",X"1A",X"6E",X"0C",
		X"F8",X"EB",X"F9",X"1D",X"15",X"12",X"10",X"00",X"10",X"00",X"00",X"F7",X"EA",X"F8",X"1C",X"14",
		X"02",X"0E",X"00",X"0E",X"00",X"0A",X"00",X"FD",X"FD",X"01",X"FD",X"12",X"06",X"00",X"06",X"00",
		X"0A",X"0F",X"FC",X"FC",X"07",X"FC",X"02",X"0E",X"00",X"0E",X"00",X"0C",X"00",X"F8",X"F8",X"01",
		X"F8",X"12",X"06",X"00",X"06",X"00",X"0C",X"0B",X"F7",X"F7",X"08",X"F7",X"04",X"1C",X"00",X"1C",
		X"00",X"00",X"00",X"E5",X"ED",X"01",X"0F",X"E4",X"1E",X"21",X"20",X"21",X"00",X"FF",X"E8",X"EC",
		X"04",X"12",X"C4",X"1E",X"79",X"26",X"4D",X"0C",X"08",X"01",X"FD",X"01",X"01",X"84",X"22",X"A5",
		X"28",X"4D",X"0A",X"09",X"01",X"FA",X"01",X"01",X"C4",X"1E",X"79",X"26",X"4D",X"0A",X"FC",X"E5",
		X"E9",X"01",X"0F",X"E4",X"22",X"21",X"24",X"21",X"00",X"FB",X"E0",X"E8",X"FC",X"0A",X"C4",X"22",
		X"79",X"28",X"4D",X"0C",X"04",X"01",X"F9",X"01",X"01",X"84",X"1E",X"A5",X"26",X"4D",X"0A",X"05",
		X"01",X"F6",X"01",X"01",X"C4",X"22",X"79",X"28",X"4D",X"0A",X"F8",X"DD",X"E5",X"F9",X"07",X"14",
		X"1E",X"00",X"1E",X"00",X"00",X"F7",X"DC",X"E4",X"F8",X"06",X"04",X"1C",X"00",X"1C",X"00",X"0C",
		X"00",X"FD",X"01",X"FD",X"FD",X"14",X"30",X"00",X"30",X"00",X"0C",X"F3",X"FC",X"EB",X"FC",X"FC",
		X"04",X"1C",X"00",X"1C",X"00",X"0A",X"00",X"01",X"01",X"F8",X"F8",X"14",X"30",X"00",X"30",X"00",
		X"0A",X"EF",X"00",X"EC",X"F7",X"F7",X"08",X"2A",X"00",X"2A",X"00",X"00",X"00",X"FB",X"E5",X"F3",
		X"01",X"E8",X"2C",X"2C",X"2E",X"2C",X"00",X"FF",X"FA",X"E8",X"F6",X"04",X"C8",X"2C",X"84",X"34",
		X"58",X"04",X"08",X"E1",X"01",X"01",X"01",X"88",X"30",X"B0",X"36",X"58",X"02",X"09",X"DE",X"01",
		X"01",X"01",X"C8",X"2C",X"84",X"34",X"58",X"02",X"FC",X"F7",X"E5",X"F3",X"01",X"E8",X"30",X"2C",
		X"32",X"2C",X"00",X"FB",X"F6",X"E0",X"EE",X"FC",X"C8",X"30",X"84",X"36",X"58",X"04",X"04",X"DD",
		X"01",X"01",X"01",X"88",X"2C",X"B0",X"34",X"58",X"02",X"05",X"DA",X"01",X"01",X"01",X"C8",X"30",
		X"84",X"36",X"58",X"02",X"F8",X"F3",X"DD",X"EB",X"F9",X"18",X"2C",X"00",X"2C",X"00",X"00",X"F7",
		X"F2",X"DC",X"EA",X"F8",X"08",X"2A",X"00",X"2A",X"00",X"04",X"00",X"01",X"FD",X"FD",X"FD",X"18",
		X"14",X"00",X"14",X"00",X"04",X"D7",X"CF",X"FC",X"FC",X"FC",X"08",X"2A",X"00",X"2A",X"00",X"02",
		X"00",X"01",X"F8",X"F8",X"F8",X"18",X"14",X"00",X"14",X"00",X"02",X"D3",X"D0",X"F7",X"F7",X"F7",
		X"C5",X"F0",X"26",X"06",X"8E",X"B7",X"14",X"3A",X"3A",X"39",X"8E",X"B7",X"32",X"30",X"02",X"58",
		X"24",X"FB",X"39",X"C5",X"F0",X"26",X"11",X"C1",X"02",X"23",X"E5",X"8E",X"B7",X"18",X"C6",X"02",
		X"30",X"02",X"5C",X"A6",X"84",X"26",X"F9",X"39",X"8E",X"B7",X"34",X"A6",X"84",X"27",X"F8",X"54",
		X"30",X"02",X"20",X"F7",X"BD",X"51",X"50",X"AE",X"84",X"2B",X"01",X"39",X"34",X"20",X"A6",X"88",
		X"51",X"27",X"52",X"EC",X"4C",X"A3",X"0C",X"2A",X"04",X"43",X"50",X"82",X"FF",X"E0",X"C8",X"54",
		X"82",X"00",X"E0",X"88",X"54",X"82",X"00",X"2A",X"3C",X"EC",X"4E",X"A3",X"0E",X"2A",X"04",X"43",
		X"50",X"82",X"FF",X"E0",X"C8",X"55",X"82",X"00",X"E0",X"88",X"55",X"82",X"00",X"2A",X"26",X"E6",
		X"02",X"E0",X"42",X"2A",X"01",X"50",X"E0",X"C8",X"56",X"E0",X"88",X"56",X"2A",X"17",X"10",X"8E",
		X"52",X"1C",X"A6",X"51",X"48",X"AB",X"51",X"48",X"AB",X"11",X"48",X"34",X"50",X"AD",X"B6",X"35",
		X"50",X"1A",X"01",X"35",X"A0",X"1C",X"FE",X"35",X"A0",X"34",X"20",X"A6",X"88",X"51",X"27",X"F5",
		X"EC",X"4C",X"A3",X"0C",X"2A",X"04",X"43",X"50",X"82",X"FF",X"E0",X"C8",X"54",X"82",X"00",X"E0",
		X"88",X"54",X"82",X"00",X"2A",X"DF",X"EC",X"4E",X"A3",X"0E",X"2A",X"04",X"43",X"50",X"82",X"FF",
		X"E0",X"C8",X"55",X"82",X"00",X"E0",X"88",X"55",X"82",X"00",X"2A",X"C9",X"C6",X"04",X"EB",X"02",
		X"E0",X"42",X"2B",X"C1",X"C1",X"10",X"22",X"BD",X"20",X"A4",X"52",X"72",X"53",X"95",X"53",X"43",
		X"52",X"78",X"52",X"75",X"52",X"72",X"53",X"95",X"52",X"72",X"53",X"43",X"52",X"78",X"52",X"75",
		X"52",X"72",X"53",X"A0",X"53",X"A0",X"52",X"72",X"52",X"73",X"52",X"73",X"52",X"72",X"53",X"AE",
		X"53",X"AE",X"52",X"73",X"52",X"73",X"52",X"73",X"52",X"72",X"52",X"76",X"52",X"76",X"52",X"73",
		X"52",X"73",X"52",X"73",X"52",X"72",X"53",X"A0",X"53",X"A0",X"52",X"74",X"52",X"74",X"52",X"74",
		X"52",X"72",X"39",X"39",X"39",X"3F",X"3F",X"39",X"C1",X"08",X"25",X"4C",X"A6",X"88",X"51",X"85",
		X"02",X"27",X"44",X"A6",X"88",X"51",X"84",X"FD",X"A7",X"88",X"51",X"26",X"19",X"A6",X"88",X"18",
		X"27",X"14",X"5F",X"A6",X"88",X"20",X"85",X"09",X"26",X"02",X"CB",X"0A",X"10",X"8E",X"02",X"46",
		X"31",X"A5",X"10",X"AF",X"88",X"29",X"CC",X"4B",X"67",X"ED",X"88",X"25",X"FC",X"EF",X"D4",X"ED",
		X"88",X"58",X"CC",X"01",X"01",X"ED",X"88",X"18",X"AE",X"88",X"22",X"EC",X"88",X"22",X"BD",X"11",
		X"1D",X"8E",X"77",X"B4",X"7E",X"E0",X"75",X"39",X"A6",X"88",X"51",X"85",X"01",X"27",X"73",X"EC",
		X"4C",X"A3",X"0C",X"2A",X"04",X"43",X"50",X"82",X"FF",X"E0",X"C8",X"54",X"82",X"00",X"C0",X"0C",
		X"82",X"00",X"2B",X"1C",X"EC",X"4E",X"A3",X"0E",X"2A",X"04",X"43",X"50",X"82",X"FF",X"E0",X"C8",
		X"55",X"82",X"00",X"C0",X"0C",X"82",X"00",X"2A",X"49",X"A6",X"88",X"51",X"85",X"01",X"27",X"42",
		X"A6",X"88",X"51",X"84",X"FE",X"A7",X"88",X"51",X"27",X"08",X"CC",X"4B",X"FF",X"ED",X"88",X"25",
		X"20",X"0A",X"A6",X"88",X"19",X"27",X"05",X"4F",X"5F",X"ED",X"88",X"2B",X"CC",X"4B",X"FE",X"ED",
		X"88",X"27",X"FC",X"EF",X"D6",X"ED",X"88",X"58",X"CC",X"01",X"01",X"ED",X"88",X"18",X"86",X"FF",
		X"A7",X"88",X"5E",X"AE",X"88",X"22",X"EC",X"88",X"20",X"BD",X"11",X"1D",X"8E",X"77",X"B7",X"7E",
		X"E0",X"75",X"39",X"7A",X"B8",X"34",X"10",X"AE",X"88",X"22",X"EC",X"2E",X"ED",X"88",X"25",X"EC",
		X"A8",X"10",X"ED",X"88",X"27",X"FC",X"EF",X"B8",X"ED",X"88",X"5A",X"FC",X"EF",X"CA",X"ED",X"88",
		X"58",X"86",X"0C",X"A7",X"88",X"5C",X"86",X"FF",X"F6",X"B7",X"48",X"27",X"13",X"CC",X"76",X"C9",
		X"ED",X"88",X"25",X"34",X"10",X"AE",X"C8",X"22",X"AE",X"88",X"1A",X"6C",X"84",X"35",X"10",X"4F",
		X"A7",X"88",X"51",X"EC",X"A8",X"22",X"BD",X"11",X"1D",X"AE",X"2C",X"B6",X"B7",X"48",X"27",X"02",
		X"AE",X"2A",X"7E",X"E0",X"75",X"0C",X"90",X"CC",X"62",X"8C",X"ED",X"14",X"6F",X"88",X"51",X"39",
		X"0C",X"90",X"10",X"AE",X"88",X"22",X"EC",X"28",X"ED",X"14",X"6F",X"88",X"51",X"39",X"A6",X"C8",
		X"51",X"81",X"02",X"26",X"0F",X"34",X"76",X"10",X"8E",X"53",X"C6",X"86",X"0D",X"C6",X"FF",X"BD",
		X"E0",X"63",X"35",X"76",X"20",X"DA",X"CC",X"0D",X"FF",X"BD",X"E0",X"66",X"86",X"96",X"A7",X"48",
		X"5F",X"6A",X"48",X"A6",X"48",X"27",X"10",X"C6",X"11",X"84",X"07",X"26",X"0A",X"5F",X"8D",X"15",
		X"86",X"04",X"BD",X"E0",X"7D",X"C6",X"11",X"8D",X"0C",X"86",X"01",X"BD",X"E0",X"7D",X"A6",X"48",
		X"26",X"DE",X"7E",X"E0",X"69",X"8E",X"1E",X"20",X"86",X"A5",X"7E",X"E0",X"25",X"10",X"AE",X"C8",
		X"22",X"E6",X"A8",X"1C",X"BD",X"51",X"63",X"EF",X"84",X"E7",X"C8",X"11",X"10",X"AE",X"C8",X"22",
		X"AE",X"24",X"AF",X"C8",X"2F",X"AE",X"26",X"AF",X"C8",X"2D",X"BD",X"69",X"26",X"20",X"11",X"10",
		X"AE",X"C8",X"22",X"AE",X"24",X"AF",X"C8",X"2F",X"AE",X"26",X"AF",X"C8",X"2D",X"BD",X"69",X"15",
		X"EC",X"A4",X"ED",X"C8",X"25",X"EC",X"22",X"ED",X"C8",X"27",X"4F",X"5F",X"ED",X"C8",X"33",X"6F",
		X"C8",X"13",X"6F",X"C8",X"57",X"6F",X"C8",X"3B",X"A6",X"A8",X"1E",X"A7",X"C8",X"51",X"BD",X"E0",
		X"B0",X"25",X"03",X"BD",X"E0",X"80",X"FC",X"EF",X"B8",X"ED",X"C8",X"5A",X"31",X"C8",X"3A",X"C6",
		X"08",X"34",X"76",X"A6",X"51",X"81",X"05",X"27",X"25",X"EE",X"C8",X"14",X"33",X"C9",X"91",X"02",
		X"96",X"9D",X"27",X"1A",X"A6",X"C8",X"BF",X"2A",X"05",X"40",X"A7",X"A4",X"20",X"10",X"E6",X"61",
		X"BD",X"E0",X"99",X"18",X"03",X"05",X"A6",X"A2",X"26",X"04",X"64",X"61",X"26",X"F0",X"35",X"F6",
		X"34",X"20",X"10",X"9E",X"66",X"8D",X"02",X"35",X"A0",X"34",X"20",X"32",X"7C",X"BD",X"E0",X"72",
		X"49",X"1F",X"89",X"BD",X"E0",X"72",X"49",X"1F",X"01",X"E6",X"64",X"3D",X"ED",X"E4",X"1F",X"10",
		X"A6",X"65",X"3D",X"ED",X"62",X"1F",X"10",X"E6",X"65",X"3D",X"E3",X"61",X"ED",X"61",X"86",X"00",
		X"A9",X"E4",X"A7",X"E4",X"1F",X"10",X"A6",X"64",X"3D",X"E3",X"61",X"ED",X"61",X"86",X"00",X"A9",
		X"E4",X"A7",X"E4",X"EC",X"E4",X"C3",X"00",X"01",X"1F",X"02",X"8E",X"91",X"02",X"A6",X"80",X"2F",
		X"FC",X"85",X"0F",X"27",X"F8",X"85",X"10",X"26",X"F4",X"31",X"3F",X"26",X"F0",X"30",X"1F",X"32",
		X"64",X"35",X"A0",X"BD",X"54",X"90",X"EC",X"81",X"27",X"1D",X"4D",X"2F",X"08",X"85",X"10",X"26",
		X"04",X"84",X"0F",X"26",X"1E",X"5D",X"2F",X"0F",X"C5",X"10",X"26",X"F9",X"C4",X"0F",X"26",X"0F",
		X"20",X"05",X"12",X"30",X"89",X"91",X"04",X"9C",X"62",X"25",X"DB",X"9E",X"60",X"20",X"D7",X"1F",
		X"98",X"30",X"01",X"A6",X"89",X"09",X"3E",X"26",X"EE",X"30",X"89",X"6E",X"FC",X"BD",X"5F",X"B1",
		X"27",X"E1",X"BD",X"5F",X"A5",X"27",X"DC",X"FC",X"B8",X"14",X"27",X"28",X"1F",X"10",X"F3",X"91",
		X"00",X"58",X"49",X"58",X"49",X"54",X"54",X"ED",X"C8",X"16",X"B0",X"B8",X"14",X"25",X"15",X"F0",
		X"B8",X"15",X"25",X"10",X"4D",X"27",X"09",X"5D",X"26",X"0A",X"81",X"03",X"23",X"B4",X"20",X"04",
		X"C1",X"03",X"23",X"AE",X"30",X"89",X"91",X"02",X"1F",X"10",X"83",X"91",X"02",X"ED",X"C8",X"14",
		X"F3",X"91",X"00",X"58",X"49",X"58",X"49",X"54",X"54",X"ED",X"C8",X"16",X"ED",X"C8",X"1C",X"ED",
		X"C8",X"1A",X"39",X"AE",X"C8",X"2F",X"6C",X"C8",X"12",X"A6",X"C8",X"12",X"46",X"24",X"02",X"30",
		X"02",X"30",X"88",X"38",X"AF",X"C8",X"29",X"BD",X"E0",X"88",X"86",X"01",X"7E",X"E0",X"7D",X"AE",
		X"C8",X"41",X"A6",X"89",X"9A",X"42",X"84",X"0F",X"27",X"08",X"A8",X"C8",X"11",X"27",X"0E",X"1A",
		X"01",X"39",X"A6",X"C8",X"11",X"AA",X"89",X"9A",X"42",X"A7",X"89",X"9A",X"42",X"1C",X"FE",X"39",
		X"6F",X"C8",X"5F",X"7C",X"B8",X"03",X"8E",X"77",X"BA",X"BD",X"E0",X"9E",X"6F",X"C8",X"39",X"6F",
		X"C8",X"13",X"FC",X"B8",X"14",X"26",X"06",X"BD",X"54",X"F3",X"EC",X"C8",X"16",X"ED",X"C8",X"16",
		X"BD",X"53",X"FD",X"6F",X"C8",X"51",X"CC",X"0C",X"0C",X"ED",X"C8",X"54",X"86",X"04",X"A7",X"C8",
		X"56",X"A6",X"42",X"8B",X"05",X"A7",X"C8",X"43",X"80",X"0C",X"A7",X"42",X"A6",X"5E",X"8B",X"0C",
		X"A7",X"5E",X"AE",X"C8",X"14",X"E6",X"89",X"91",X"02",X"54",X"54",X"C4",X"3C",X"CB",X"02",X"E7",
		X"C8",X"5E",X"6F",X"C8",X"51",X"FC",X"EF",X"C0",X"ED",X"C8",X"5A",X"6F",X"C8",X"40",X"86",X"0F",
		X"A7",X"C8",X"44",X"EC",X"C8",X"14",X"AE",X"C8",X"16",X"34",X"16",X"AE",X"C8",X"41",X"96",X"68",
		X"2A",X"06",X"BD",X"54",X"F3",X"AE",X"C8",X"14",X"AF",X"C8",X"41",X"A6",X"C8",X"11",X"AA",X"89",
		X"9A",X"42",X"A7",X"89",X"9A",X"42",X"1F",X"10",X"F3",X"91",X"00",X"58",X"49",X"58",X"49",X"54",
		X"54",X"ED",X"C8",X"3E",X"35",X"16",X"ED",X"C8",X"14",X"AF",X"C8",X"16",X"AF",X"C8",X"1C",X"AF",
		X"C8",X"1A",X"BD",X"55",X"83",X"BD",X"55",X"9F",X"E6",X"C8",X"43",X"E1",X"42",X"27",X"12",X"2D",
		X"09",X"6A",X"5E",X"6C",X"C8",X"5E",X"6C",X"42",X"20",X"07",X"6C",X"5E",X"6A",X"C8",X"5E",X"6A",
		X"42",X"EC",X"C8",X"3E",X"10",X"A3",X"C8",X"16",X"27",X"78",X"6D",X"C8",X"40",X"2B",X"18",X"2E",
		X"37",X"A0",X"C8",X"16",X"24",X"01",X"40",X"E0",X"C8",X"17",X"24",X"01",X"50",X"34",X"02",X"E0",
		X"E0",X"12",X"E7",X"C8",X"40",X"2E",X"21",X"A6",X"C8",X"16",X"A1",X"C8",X"3E",X"26",X"05",X"6F",
		X"C8",X"40",X"20",X"14",X"25",X"05",X"8E",X"65",X"00",X"20",X"03",X"8E",X"65",X"0B",X"BD",X"72",
		X"96",X"63",X"C8",X"13",X"2B",X"9C",X"20",X"21",X"E6",X"C8",X"17",X"E1",X"C8",X"3F",X"26",X"05",
		X"6F",X"C8",X"40",X"20",X"8D",X"25",X"05",X"8E",X"64",X"F5",X"20",X"03",X"8E",X"65",X"16",X"BD",
		X"72",X"96",X"63",X"C8",X"13",X"10",X"2B",X"FF",X"79",X"EC",X"04",X"E3",X"C8",X"14",X"ED",X"C8",
		X"14",X"EC",X"06",X"E3",X"C8",X"16",X"ED",X"C8",X"16",X"ED",X"C8",X"1C",X"ED",X"C8",X"1A",X"7E",
		X"56",X"62",X"A6",X"C8",X"44",X"A7",X"C8",X"40",X"27",X"12",X"64",X"C8",X"44",X"BD",X"55",X"83",
		X"BD",X"55",X"9F",X"10",X"25",X"FF",X"0C",X"6A",X"C8",X"40",X"26",X"F1",X"BD",X"55",X"83",X"BD",
		X"55",X"9F",X"10",X"25",X"FE",X"FD",X"BD",X"55",X"83",X"BD",X"55",X"9F",X"10",X"25",X"FE",X"F3",
		X"AE",X"C8",X"14",X"E6",X"89",X"91",X"02",X"54",X"54",X"C4",X"3C",X"A6",X"42",X"80",X"05",X"34",
		X"02",X"E1",X"E0",X"27",X"14",X"2D",X"09",X"6A",X"5E",X"6C",X"C8",X"5E",X"6C",X"42",X"20",X"CC",
		X"6C",X"5E",X"6A",X"C8",X"5E",X"6A",X"42",X"20",X"C3",X"BD",X"55",X"83",X"BD",X"55",X"9F",X"10",
		X"25",X"FE",X"C0",X"8E",X"77",X"C0",X"BD",X"E0",X"75",X"7A",X"B8",X"03",X"26",X"06",X"8E",X"77",
		X"BD",X"BD",X"E0",X"9E",X"6F",X"C8",X"3F",X"6F",X"C8",X"42",X"6F",X"C8",X"45",X"6F",X"C8",X"48",
		X"86",X"10",X"A7",X"C8",X"12",X"BD",X"54",X"0C",X"6F",X"43",X"6F",X"C8",X"20",X"86",X"04",X"8E",
		X"50",X"1C",X"E6",X"C8",X"16",X"E1",X"C8",X"17",X"25",X"05",X"86",X"08",X"8E",X"50",X"B6",X"A7",
		X"C8",X"10",X"A7",X"C8",X"21",X"AF",X"C8",X"1E",X"AE",X"C8",X"14",X"A6",X"89",X"91",X"02",X"A7",
		X"C8",X"24",X"A6",X"89",X"9A",X"42",X"AA",X"C8",X"11",X"A7",X"89",X"9A",X"42",X"6F",X"C8",X"3E",
		X"CC",X"0C",X"0C",X"ED",X"C8",X"54",X"86",X"08",X"A7",X"C8",X"56",X"4F",X"5F",X"ED",X"4A",X"6F",
		X"C8",X"3D",X"CC",X"6F",X"1D",X"ED",X"C8",X"27",X"CC",X"72",X"D6",X"ED",X"C8",X"25",X"FC",X"EF",
		X"E8",X"ED",X"C8",X"5A",X"7C",X"B8",X"33",X"7E",X"58",X"27",X"E6",X"24",X"6C",X"C8",X"13",X"3A",
		X"BD",X"72",X"96",X"AE",X"C8",X"2F",X"E6",X"23",X"3A",X"AF",X"C8",X"29",X"A6",X"C8",X"51",X"2A",
		X"03",X"BD",X"59",X"91",X"BD",X"59",X"91",X"BD",X"59",X"91",X"10",X"AE",X"C8",X"1E",X"A6",X"A4",
		X"48",X"2A",X"0F",X"AE",X"C8",X"14",X"A6",X"C8",X"11",X"43",X"A4",X"89",X"9A",X"42",X"A7",X"89",
		X"9A",X"42",X"8E",X"64",X"EA",X"20",X"0B",X"10",X"AE",X"C8",X"1E",X"8E",X"64",X"EA",X"A6",X"A4",
		X"2B",X"B8",X"E6",X"22",X"6F",X"C8",X"13",X"3A",X"BD",X"5F",X"CE",X"24",X"07",X"A6",X"C8",X"51",
		X"10",X"2B",X"09",X"AB",X"A6",X"43",X"27",X"44",X"BD",X"72",X"96",X"A6",X"A4",X"48",X"2A",X"3C",
		X"EC",X"04",X"E3",X"C8",X"14",X"ED",X"C8",X"14",X"EC",X"06",X"E3",X"C8",X"16",X"ED",X"C8",X"16",
		X"ED",X"C8",X"1C",X"ED",X"C8",X"1A",X"AE",X"C8",X"14",X"A6",X"89",X"90",X"C1",X"2A",X"08",X"81",
		X"81",X"27",X"04",X"40",X"A7",X"C8",X"3A",X"A6",X"C8",X"51",X"2B",X"09",X"A6",X"89",X"91",X"02",
		X"BD",X"59",X"47",X"20",X"07",X"BD",X"59",X"1E",X"10",X"25",X"09",X"63",X"A6",X"A4",X"85",X"10",
		X"26",X"07",X"AD",X"D8",X"25",X"10",X"AE",X"C8",X"1E",X"A6",X"43",X"8E",X"64",X"B4",X"E6",X"86",
		X"86",X"0B",X"E6",X"A5",X"3D",X"2A",X"02",X"80",X"0B",X"31",X"AB",X"E6",X"22",X"8E",X"64",X"EA",
		X"3A",X"EC",X"04",X"E3",X"C8",X"14",X"1F",X"01",X"A6",X"A4",X"48",X"2A",X"36",X"E6",X"89",X"9A",
		X"42",X"27",X"26",X"A6",X"C8",X"51",X"2A",X"19",X"C4",X"0F",X"27",X"15",X"C1",X"02",X"22",X"11",
		X"BD",X"51",X"50",X"AE",X"84",X"2A",X"0A",X"1E",X"13",X"BD",X"5F",X"31",X"1E",X"13",X"6E",X"D8",
		X"F4",X"10",X"AE",X"C8",X"1E",X"6F",X"43",X"20",X"B0",X"AF",X"C8",X"31",X"EA",X"C8",X"11",X"E7",
		X"89",X"9A",X"42",X"A6",X"A4",X"85",X"20",X"27",X"0A",X"A6",X"89",X"91",X"02",X"85",X"10",X"27",
		X"02",X"31",X"2B",X"10",X"AF",X"C8",X"1E",X"AE",X"C8",X"2F",X"E6",X"21",X"3A",X"AF",X"C8",X"29",
		X"A6",X"C8",X"51",X"2A",X"02",X"8D",X"7A",X"8D",X"78",X"8D",X"76",X"7E",X"58",X"27",X"A6",X"89",
		X"91",X"02",X"85",X"0F",X"27",X"0F",X"BC",X"B7",X"40",X"26",X"0D",X"7D",X"B7",X"43",X"27",X"35",
		X"B6",X"B7",X"42",X"20",X"30",X"1A",X"01",X"39",X"BC",X"B7",X"44",X"26",X"0A",X"7D",X"B7",X"47",
		X"27",X"23",X"B6",X"B7",X"46",X"20",X"1E",X"BC",X"B7",X"49",X"27",X"1E",X"BC",X"B7",X"50",X"27",
		X"1E",X"BC",X"B7",X"57",X"27",X"1E",X"BC",X"B7",X"5E",X"27",X"1E",X"BC",X"B7",X"65",X"27",X"1E",
		X"BC",X"B7",X"6C",X"27",X"1E",X"A7",X"C8",X"24",X"5F",X"39",X"B6",X"B7",X"4B",X"20",X"17",X"B6",
		X"B7",X"52",X"20",X"12",X"B6",X"B7",X"59",X"20",X"0D",X"B6",X"B7",X"60",X"20",X"08",X"B6",X"B7",
		X"67",X"20",X"03",X"B6",X"B7",X"6E",X"A7",X"C8",X"24",X"E6",X"C8",X"3D",X"27",X"D7",X"1C",X"FE",
		X"39",X"A6",X"C8",X"51",X"26",X"07",X"A6",X"C8",X"5C",X"10",X"27",X"08",X"7B",X"AD",X"D8",X"27",
		X"8E",X"64",X"BD",X"A6",X"C8",X"21",X"26",X"03",X"A6",X"C8",X"10",X"A7",X"C8",X"10",X"E6",X"86",
		X"AE",X"C8",X"2D",X"3A",X"AF",X"C8",X"2B",X"BD",X"E0",X"88",X"86",X"01",X"7E",X"E0",X"7D",X"10",
		X"AE",X"C8",X"22",X"C6",X"01",X"A6",X"51",X"81",X"02",X"26",X"02",X"C6",X"02",X"E7",X"C8",X"20",
		X"E7",X"C8",X"10",X"6F",X"C8",X"21",X"9E",X"25",X"A6",X"A8",X"1D",X"30",X"86",X"86",X"05",X"BD",
		X"E0",X"83",X"ED",X"C8",X"16",X"ED",X"C8",X"1C",X"ED",X"C8",X"1A",X"86",X"08",X"A7",X"C8",X"56",
		X"BD",X"E0",X"B0",X"25",X"03",X"BD",X"E0",X"80",X"EE",X"C8",X"44",X"2B",X"F3",X"DE",X"21",X"BD",
		X"53",X"FD",X"96",X"68",X"2B",X"09",X"FC",X"E0",X"8E",X"ED",X"C8",X"25",X"ED",X"C8",X"27",X"FC",
		X"EF",X"BA",X"ED",X"C8",X"5A",X"6F",X"43",X"A6",X"C8",X"20",X"48",X"8E",X"5A",X"54",X"EC",X"86",
		X"ED",X"C8",X"1E",X"AE",X"C8",X"14",X"A6",X"89",X"91",X"02",X"A7",X"C8",X"24",X"6F",X"C8",X"3E",
		X"6F",X"C8",X"3B",X"6F",X"C8",X"12",X"CC",X"0C",X"0C",X"ED",X"C8",X"54",X"86",X"08",X"A7",X"C8",
		X"56",X"CC",X"00",X"00",X"ED",X"4A",X"10",X"AE",X"C8",X"1E",X"AE",X"C8",X"2F",X"E6",X"21",X"3A",
		X"AF",X"C8",X"29",X"39",X"4E",X"E8",X"4E",X"E8",X"4F",X"82",X"00",X"00",X"50",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"B6",X"1F",X"89",X"BD",X"51",X"50",X"AE",X"84",X"A6",X"11",X"81",
		X"03",X"26",X"15",X"A6",X"88",X"51",X"2F",X"07",X"34",X"10",X"BD",X"53",X"43",X"35",X"10",X"A6",
		X"88",X"51",X"2A",X"03",X"BD",X"5F",X"31",X"39",X"81",X"04",X"26",X"0B",X"34",X"10",X"BD",X"52",
		X"7C",X"35",X"10",X"BD",X"52",X"F9",X"39",X"3F",X"39",X"34",X"30",X"6F",X"C8",X"3D",X"10",X"AE",
		X"C8",X"22",X"AE",X"A8",X"14",X"2A",X"04",X"6F",X"07",X"6C",X"04",X"35",X"B0",X"BD",X"59",X"BF",
		X"BD",X"5A",X"99",X"6F",X"C8",X"51",X"6F",X"C8",X"5F",X"6F",X"C8",X"20",X"6F",X"C8",X"48",X"FC",
		X"E0",X"8E",X"ED",X"C8",X"5A",X"86",X"0A",X"A7",X"C8",X"37",X"AE",X"C8",X"14",X"A6",X"89",X"9A",
		X"42",X"27",X"2E",X"6A",X"C8",X"37",X"26",X"1E",X"85",X"0F",X"27",X"02",X"84",X"0F",X"81",X"02",
		X"22",X"1C",X"10",X"8E",X"31",X"28",X"A6",X"51",X"81",X"02",X"27",X"04",X"10",X"8E",X"31",X"4C",
		X"BD",X"59",X"C3",X"7E",X"5A",X"B3",X"8E",X"5A",X"CA",X"86",X"02",X"7E",X"E0",X"6C",X"BD",X"5A",
		X"66",X"96",X"90",X"27",X"10",X"8E",X"77",X"48",X"A6",X"C8",X"11",X"81",X"01",X"27",X"03",X"8E",
		X"77",X"4B",X"BD",X"E0",X"9E",X"A6",X"C8",X"11",X"AE",X"C8",X"14",X"A7",X"89",X"9A",X"42",X"AE",
		X"C8",X"22",X"A6",X"88",X"1F",X"A7",X"C8",X"37",X"FC",X"EF",X"CE",X"ED",X"C8",X"5A",X"6F",X"C8",
		X"51",X"6F",X"C8",X"35",X"6F",X"C8",X"39",X"AD",X"D8",X"25",X"A6",X"43",X"A7",X"C8",X"34",X"20",
		X"03",X"AD",X"D8",X"25",X"A6",X"43",X"27",X"05",X"A1",X"C8",X"34",X"26",X"29",X"A7",X"C8",X"34",
		X"A6",X"C8",X"35",X"27",X"0E",X"AD",X"D8",X"25",X"BD",X"5F",X"74",X"6C",X"C8",X"39",X"BD",X"5F",
		X"74",X"20",X"09",X"BD",X"5F",X"81",X"6C",X"C8",X"39",X"BD",X"5F",X"81",X"6C",X"C8",X"39",X"A6",
		X"C8",X"39",X"81",X"B4",X"25",X"CB",X"8E",X"77",X"4E",X"A6",X"C8",X"11",X"81",X"01",X"27",X"03",
		X"8E",X"77",X"51",X"BD",X"E0",X"9E",X"FC",X"EF",X"BA",X"ED",X"C8",X"5A",X"6F",X"C8",X"20",X"86",
		X"01",X"A7",X"C8",X"51",X"E6",X"C8",X"11",X"BD",X"51",X"63",X"EF",X"84",X"7E",X"5B",X"D4",X"E6",
		X"24",X"6C",X"C8",X"13",X"3A",X"BD",X"72",X"96",X"AE",X"C8",X"2F",X"E6",X"23",X"3A",X"AF",X"C8",
		X"29",X"BD",X"5F",X"74",X"BD",X"5F",X"74",X"10",X"AE",X"C8",X"1E",X"A6",X"A4",X"48",X"2A",X"0F",
		X"AE",X"C8",X"14",X"A6",X"C8",X"11",X"43",X"A4",X"89",X"9A",X"42",X"A7",X"89",X"9A",X"42",X"8E",
		X"64",X"EA",X"20",X"0B",X"10",X"AE",X"C8",X"1E",X"8E",X"64",X"EA",X"A6",X"A4",X"2B",X"C0",X"E6",
		X"22",X"6F",X"C8",X"13",X"3A",X"B6",X"B8",X"14",X"26",X"15",X"EC",X"C8",X"16",X"B1",X"B8",X"29",
		X"23",X"05",X"F1",X"B8",X"29",X"22",X"08",X"0C",X"90",X"6F",X"C8",X"51",X"7E",X"62",X"97",X"BD",
		X"5F",X"CE",X"24",X"12",X"96",X"90",X"27",X"0E",X"A6",X"51",X"40",X"97",X"90",X"CC",X"00",X"F0",
		X"BD",X"E0",X"66",X"7E",X"E0",X"69",X"A6",X"43",X"27",X"2F",X"BD",X"72",X"96",X"A6",X"A4",X"48",
		X"2A",X"34",X"EC",X"04",X"E3",X"C8",X"14",X"ED",X"C8",X"14",X"EC",X"06",X"E3",X"C8",X"16",X"ED",
		X"C8",X"16",X"ED",X"C8",X"1C",X"ED",X"C8",X"1A",X"AE",X"C8",X"14",X"A6",X"89",X"90",X"C1",X"2A",
		X"08",X"81",X"81",X"27",X"04",X"40",X"A7",X"C8",X"3A",X"AE",X"C8",X"14",X"BD",X"59",X"1E",X"25",
		X"B7",X"27",X"03",X"BD",X"5E",X"A6",X"AD",X"D8",X"25",X"10",X"AE",X"C8",X"1E",X"A6",X"43",X"8E",
		X"64",X"B4",X"E6",X"86",X"86",X"0B",X"E6",X"A5",X"3D",X"2A",X"02",X"80",X"0B",X"31",X"AB",X"E6",
		X"22",X"8E",X"64",X"EA",X"3A",X"EC",X"04",X"E3",X"C8",X"14",X"1F",X"01",X"A6",X"A4",X"48",X"10",
		X"2A",X"00",X"5C",X"E6",X"89",X"9A",X"42",X"27",X"47",X"C4",X"0F",X"27",X"3A",X"E1",X"C8",X"11",
		X"27",X"3E",X"C1",X"02",X"23",X"31",X"34",X"10",X"BD",X"51",X"50",X"AE",X"84",X"2A",X"26",X"A6",
		X"88",X"51",X"2E",X"21",X"27",X"11",X"BD",X"5F",X"31",X"35",X"10",X"E6",X"89",X"9A",X"42",X"C4",
		X"F0",X"E7",X"89",X"9A",X"42",X"20",X"19",X"35",X"10",X"E6",X"89",X"9A",X"42",X"C4",X"F0",X"E7",
		X"89",X"9A",X"42",X"20",X"0B",X"35",X"10",X"10",X"AE",X"C8",X"1E",X"6F",X"43",X"7E",X"5C",X"5D",
		X"AF",X"C8",X"31",X"EA",X"C8",X"11",X"E7",X"89",X"9A",X"42",X"BD",X"5F",X"A5",X"27",X"2B",X"A6",
		X"A4",X"85",X"20",X"27",X"0A",X"A6",X"89",X"91",X"02",X"85",X"10",X"27",X"02",X"31",X"2B",X"10",
		X"AF",X"C8",X"1E",X"E6",X"25",X"E7",X"C8",X"48",X"AE",X"C8",X"2F",X"E6",X"21",X"3A",X"AF",X"C8",
		X"29",X"BD",X"5F",X"74",X"BD",X"5F",X"74",X"7E",X"5B",X"D4",X"34",X"10",X"10",X"AF",X"C8",X"1E",
		X"E6",X"25",X"E7",X"C8",X"48",X"AE",X"C8",X"2F",X"E6",X"21",X"3A",X"AF",X"C8",X"29",X"35",X"10",
		X"BD",X"5E",X"67",X"A6",X"22",X"34",X"02",X"1F",X"10",X"F3",X"91",X"00",X"58",X"49",X"58",X"49",
		X"54",X"54",X"1E",X"89",X"ED",X"C8",X"16",X"58",X"58",X"44",X"56",X"44",X"56",X"B3",X"91",X"00",
		X"1F",X"01",X"BD",X"5E",X"67",X"86",X"11",X"A7",X"25",X"10",X"AF",X"C8",X"40",X"C6",X"04",X"A6",
		X"22",X"A0",X"E0",X"46",X"2A",X"02",X"40",X"50",X"44",X"A7",X"C8",X"33",X"A7",X"C8",X"34",X"E7",
		X"C8",X"36",X"A6",X"89",X"9A",X"42",X"27",X"07",X"34",X"10",X"BD",X"5A",X"66",X"35",X"10",X"A6",
		X"C8",X"11",X"A7",X"89",X"9A",X"42",X"AE",X"C8",X"14",X"A6",X"89",X"9A",X"42",X"84",X"0F",X"A1",
		X"C8",X"11",X"26",X"08",X"A8",X"89",X"9A",X"42",X"A7",X"89",X"9A",X"42",X"AE",X"C8",X"31",X"A6",
		X"89",X"9A",X"42",X"84",X"0F",X"A1",X"C8",X"11",X"26",X"08",X"A8",X"89",X"9A",X"42",X"A7",X"89",
		X"9A",X"42",X"E6",X"C8",X"11",X"BD",X"51",X"50",X"4F",X"5F",X"ED",X"84",X"6F",X"C8",X"51",X"6F",
		X"C8",X"35",X"BD",X"E0",X"88",X"86",X"01",X"BD",X"E0",X"7D",X"BD",X"E0",X"88",X"86",X"01",X"BD",
		X"E0",X"7D",X"10",X"AE",X"C8",X"1E",X"8E",X"64",X"EA",X"E6",X"24",X"3A",X"BD",X"72",X"96",X"AE",
		X"C8",X"2F",X"E6",X"23",X"3A",X"AF",X"C8",X"29",X"BD",X"E0",X"88",X"86",X"01",X"BD",X"E0",X"7D",
		X"BD",X"E0",X"88",X"86",X"01",X"BD",X"E0",X"7D",X"10",X"AE",X"C8",X"1E",X"8E",X"64",X"EA",X"E6",
		X"24",X"3A",X"BD",X"72",X"96",X"7C",X"B8",X"01",X"8E",X"77",X"69",X"BD",X"E0",X"9E",X"8E",X"77",
		X"6F",X"BD",X"E0",X"75",X"FC",X"E0",X"8E",X"ED",X"C8",X"58",X"6F",X"C8",X"5E",X"FC",X"EF",X"C4",
		X"ED",X"C8",X"5A",X"BD",X"5E",X"84",X"6A",X"C8",X"5E",X"A6",X"C8",X"5E",X"81",X"F0",X"26",X"F3",
		X"BD",X"5E",X"7C",X"6A",X"5E",X"6C",X"C8",X"35",X"6A",X"C8",X"33",X"26",X"F3",X"BD",X"5E",X"7C",
		X"6C",X"5E",X"6A",X"C8",X"35",X"6A",X"C8",X"34",X"26",X"F3",X"8E",X"77",X"72",X"BD",X"E0",X"75",
		X"BD",X"5E",X"84",X"6C",X"C8",X"5E",X"26",X"F8",X"AE",X"C8",X"40",X"6F",X"05",X"EC",X"C8",X"16",
		X"BD",X"59",X"E2",X"7A",X"B8",X"01",X"2E",X"0C",X"8E",X"77",X"6C",X"BD",X"E0",X"9E",X"8E",X"77",
		X"75",X"BD",X"E0",X"75",X"7E",X"5B",X"86",X"10",X"8E",X"B7",X"83",X"31",X"26",X"AC",X"A4",X"26",
		X"FA",X"4F",X"5F",X"ED",X"A4",X"A7",X"25",X"6F",X"89",X"90",X"C1",X"39",X"E6",X"C8",X"36",X"1D",
		X"E3",X"5A",X"ED",X"5A",X"AE",X"C8",X"2F",X"6C",X"C8",X"12",X"A6",X"C8",X"12",X"81",X"03",X"25",
		X"04",X"4F",X"A7",X"C8",X"12",X"48",X"30",X"86",X"30",X"88",X"38",X"AF",X"C8",X"29",X"BD",X"E0",
		X"88",X"86",X"01",X"7E",X"E0",X"7D",X"34",X"36",X"10",X"AE",X"C8",X"14",X"8E",X"B7",X"42",X"30",
		X"07",X"10",X"AC",X"84",X"26",X"F9",X"EC",X"03",X"27",X"75",X"34",X"16",X"10",X"8E",X"60",X"56",
		X"86",X"0F",X"C6",X"FF",X"BD",X"E0",X"63",X"35",X"16",X"25",X"64",X"10",X"BF",X"B7",X"76",X"AF",
		X"A8",X"37",X"7F",X"B7",X"74",X"F3",X"91",X"00",X"58",X"49",X"58",X"49",X"54",X"54",X"ED",X"A8",
		X"16",X"ED",X"A8",X"1C",X"ED",X"A8",X"1A",X"A6",X"C8",X"36",X"A7",X"A8",X"36",X"6F",X"A8",X"51",
		X"4F",X"5F",X"ED",X"03",X"10",X"AE",X"05",X"6A",X"A4",X"86",X"00",X"A7",X"3F",X"FC",X"EF",X"CC",
		X"ED",X"C8",X"58",X"86",X"11",X"A7",X"C8",X"5D",X"6A",X"C8",X"3D",X"AE",X"C8",X"22",X"AE",X"88",
		X"14",X"A6",X"07",X"8B",X"99",X"19",X"A7",X"07",X"6C",X"04",X"CC",X"15",X"02",X"BD",X"11",X"1D",
		X"8E",X"77",X"57",X"BD",X"E0",X"75",X"8E",X"78",X"07",X"BD",X"E0",X"9E",X"7C",X"B7",X"73",X"35",
		X"B6",X"34",X"30",X"6C",X"C8",X"3D",X"10",X"AE",X"C8",X"22",X"10",X"AE",X"A8",X"14",X"A6",X"27",
		X"8B",X"01",X"19",X"A7",X"27",X"6C",X"24",X"6F",X"88",X"51",X"FC",X"EF",X"CC",X"ED",X"C8",X"58",
		X"34",X"10",X"AE",X"88",X"22",X"A6",X"88",X"1F",X"A7",X"C8",X"5D",X"EC",X"88",X"20",X"BD",X"11",
		X"1D",X"8E",X"77",X"E1",X"BD",X"E0",X"75",X"AE",X"E4",X"AE",X"88",X"22",X"EC",X"08",X"35",X"10",
		X"ED",X"14",X"35",X"B0",X"A6",X"C8",X"12",X"34",X"02",X"AD",X"D8",X"27",X"35",X"02",X"BD",X"66",
		X"37",X"5F",X"A6",X"C8",X"21",X"26",X"0A",X"A6",X"C8",X"10",X"6D",X"C8",X"3B",X"26",X"02",X"C6",
		X"08",X"8E",X"64",X"BD",X"EB",X"86",X"AE",X"C8",X"2D",X"3A",X"AF",X"C8",X"2B",X"BD",X"E0",X"88",
		X"86",X"01",X"7E",X"E0",X"7D",X"A6",X"89",X"90",X"C1",X"2A",X"03",X"81",X"81",X"39",X"1C",X"FB",
		X"39",X"BC",X"B7",X"4C",X"27",X"17",X"BC",X"B7",X"53",X"27",X"12",X"BC",X"B7",X"5A",X"27",X"0D",
		X"BC",X"B7",X"61",X"27",X"08",X"BC",X"B7",X"68",X"27",X"03",X"BC",X"B7",X"6F",X"39",X"B6",X"B8",
		X"1A",X"A1",X"42",X"26",X"42",X"EC",X"C8",X"16",X"F0",X"B8",X"15",X"2A",X"01",X"50",X"B0",X"B8",
		X"14",X"2A",X"01",X"40",X"34",X"02",X"E1",X"E0",X"27",X"1E",X"2E",X"0F",X"7D",X"B7",X"3C",X"27",
		X"05",X"B1",X"B7",X"3C",X"22",X"12",X"B7",X"B7",X"3C",X"20",X"0D",X"7D",X"B7",X"3D",X"27",X"05",
		X"F1",X"B7",X"3D",X"22",X"03",X"F7",X"B7",X"3D",X"81",X"01",X"22",X"09",X"C1",X"01",X"22",X"05",
		X"8D",X"08",X"1A",X"01",X"39",X"8D",X"03",X"1C",X"FE",X"39",X"6D",X"C8",X"51",X"2A",X"14",X"34",
		X"02",X"E1",X"E0",X"27",X"1C",X"22",X"0D",X"34",X"04",X"AB",X"E0",X"B1",X"B7",X"3F",X"22",X"03",
		X"B7",X"B7",X"3F",X"39",X"34",X"02",X"EB",X"E0",X"F1",X"B7",X"3E",X"22",X"03",X"F7",X"B7",X"3E",
		X"39",X"34",X"04",X"AB",X"E0",X"B1",X"B7",X"3F",X"22",X"03",X"B7",X"B7",X"3F",X"B1",X"B7",X"3E",
		X"22",X"03",X"B7",X"B7",X"3E",X"39",X"CC",X"32",X"24",X"ED",X"C8",X"22",X"6F",X"C8",X"11",X"BD",
		X"54",X"0C",X"FC",X"EF",X"C2",X"ED",X"C8",X"5A",X"6F",X"43",X"6F",X"C8",X"20",X"86",X"04",X"AE",
		X"5A",X"8C",X"00",X"8B",X"25",X"02",X"86",X"08",X"A7",X"43",X"6F",X"C8",X"3E",X"CC",X"0C",X"0C",
		X"ED",X"C8",X"54",X"86",X"08",X"A7",X"C8",X"56",X"CC",X"00",X"00",X"ED",X"4A",X"E6",X"C8",X"3E",
		X"8E",X"61",X"14",X"E6",X"85",X"8E",X"03",X"12",X"A6",X"43",X"81",X"04",X"27",X"02",X"30",X"08",
		X"6A",X"5E",X"5A",X"58",X"3A",X"AF",X"C8",X"29",X"6C",X"C8",X"3E",X"E6",X"C8",X"3E",X"C1",X"1E",
		X"24",X"0B",X"BD",X"E0",X"88",X"8E",X"60",X"8D",X"86",X"01",X"7E",X"E0",X"6C",X"86",X"05",X"A7",
		X"C8",X"12",X"A7",X"C8",X"3E",X"AE",X"C8",X"37",X"4F",X"5F",X"ED",X"84",X"A7",X"02",X"11",X"B3",
		X"B7",X"76",X"26",X"03",X"FF",X"B7",X"74",X"BD",X"61",X"32",X"10",X"25",X"00",X"F6",X"A6",X"5E",
		X"81",X"C0",X"25",X"05",X"8E",X"61",X"03",X"20",X"07",X"81",X"10",X"22",X"0C",X"8E",X"61",X"0B",
		X"E6",X"43",X"E6",X"85",X"E7",X"43",X"E7",X"C8",X"20",X"BD",X"E0",X"88",X"8E",X"60",X"D7",X"86",
		X"02",X"7E",X"E0",X"6C",X"01",X"02",X"00",X"01",X"00",X"00",X"00",X"02",X"04",X"08",X"00",X"04",
		X"00",X"00",X"00",X"08",X"01",X"02",X"02",X"03",X"03",X"03",X"03",X"03",X"03",X"02",X"02",X"02",
		X"01",X"01",X"01",X"01",X"02",X"02",X"03",X"03",X"03",X"03",X"03",X"03",X"02",X"02",X"04",X"04",
		X"04",X"04",X"E6",X"43",X"BD",X"72",X"8D",X"A6",X"C8",X"13",X"88",X"01",X"A7",X"C8",X"13",X"26",
		X"36",X"EC",X"04",X"E3",X"C8",X"14",X"ED",X"C8",X"14",X"EC",X"06",X"E3",X"C8",X"16",X"ED",X"C8",
		X"16",X"10",X"8E",X"61",X"B6",X"A6",X"43",X"85",X"09",X"26",X"04",X"10",X"8E",X"61",X"C5",X"EC",
		X"A1",X"81",X"80",X"27",X"12",X"E3",X"C8",X"14",X"1F",X"01",X"A6",X"89",X"91",X"02",X"2A",X"EF",
		X"81",X"81",X"27",X"EB",X"A7",X"C8",X"3A",X"6A",X"C8",X"12",X"2E",X"23",X"86",X"05",X"A7",X"C8",
		X"12",X"A6",X"C8",X"3E",X"8B",X"02",X"81",X"02",X"23",X"01",X"4F",X"A7",X"C8",X"3E",X"8E",X"61",
		X"AD",X"E6",X"43",X"E6",X"85",X"EB",X"C8",X"3E",X"8E",X"03",X"02",X"3A",X"AF",X"C8",X"29",X"EC",
		X"5A",X"2B",X"08",X"83",X"01",X"2C",X"24",X"03",X"1C",X"FE",X"39",X"1A",X"01",X"39",X"00",X"04",
		X"00",X"08",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"40",X"FF",X"C0",X"00",X"80",X"FF",X"80",
		X"00",X"C0",X"FF",X"40",X"80",X"00",X"00",X"00",X"01",X"FF",X"FF",X"00",X"02",X"FF",X"FE",X"00",
		X"03",X"FF",X"FD",X"80",X"11",X"B3",X"B7",X"74",X"26",X"03",X"7F",X"B7",X"74",X"7A",X"B7",X"73",
		X"26",X"06",X"8E",X"78",X"0A",X"BD",X"E0",X"9E",X"6F",X"5D",X"6F",X"5E",X"7E",X"E0",X"69",X"8E",
		X"77",X"ED",X"BD",X"E0",X"75",X"AE",X"C8",X"22",X"8D",X"4D",X"AE",X"C8",X"22",X"30",X"88",X"24",
		X"8C",X"31",X"B8",X"22",X"10",X"AF",X"C8",X"22",X"0C",X"90",X"86",X"01",X"BD",X"E0",X"7D",X"7C",
		X"B8",X"34",X"7E",X"55",X"C0",X"7E",X"E0",X"69",X"8D",X"2D",X"B6",X"B7",X"48",X"26",X"25",X"FC",
		X"EF",X"C2",X"ED",X"C8",X"5A",X"8E",X"03",X"26",X"AF",X"C8",X"29",X"CC",X"FF",X"1E",X"A7",X"48",
		X"E7",X"C8",X"39",X"86",X"01",X"BD",X"E0",X"7D",X"EC",X"5E",X"83",X"00",X"80",X"ED",X"5E",X"6A",
		X"C8",X"39",X"26",X"EF",X"7E",X"E0",X"69",X"A6",X"C8",X"5F",X"27",X"06",X"6F",X"C8",X"5F",X"7A",
		X"B8",X"26",X"0A",X"90",X"AE",X"C8",X"14",X"A6",X"89",X"9A",X"42",X"84",X"0F",X"A1",X"C8",X"11",
		X"26",X"08",X"A8",X"89",X"9A",X"42",X"A7",X"89",X"9A",X"42",X"AE",X"C8",X"31",X"A6",X"89",X"9A",
		X"42",X"84",X"0F",X"A1",X"C8",X"11",X"26",X"08",X"A8",X"89",X"9A",X"42",X"A7",X"89",X"9A",X"42",
		X"E6",X"C8",X"11",X"BD",X"51",X"50",X"CC",X"00",X"00",X"ED",X"84",X"39",X"6F",X"C8",X"5E",X"8E",
		X"77",X"66",X"BD",X"E0",X"75",X"20",X"0E",X"86",X"01",X"A7",X"C8",X"5E",X"8E",X"77",X"63",X"BD",
		X"E0",X"75",X"7C",X"B8",X"21",X"A6",X"51",X"BD",X"68",X"3F",X"AE",X"C8",X"14",X"A6",X"89",X"9A",
		X"42",X"84",X"0F",X"A1",X"C8",X"11",X"26",X"08",X"A8",X"89",X"9A",X"42",X"A7",X"89",X"9A",X"42",
		X"AE",X"C8",X"31",X"A6",X"89",X"9A",X"42",X"84",X"0F",X"A1",X"C8",X"11",X"26",X"08",X"A8",X"89",
		X"9A",X"42",X"A7",X"89",X"9A",X"42",X"4F",X"E6",X"C8",X"11",X"BD",X"51",X"50",X"CC",X"00",X"00",
		X"ED",X"84",X"FC",X"E0",X"8E",X"ED",X"C8",X"58",X"FC",X"EF",X"E6",X"6D",X"C8",X"5E",X"27",X"03",
		X"FC",X"EF",X"C8",X"ED",X"C8",X"5A",X"BD",X"E0",X"88",X"86",X"01",X"BD",X"E0",X"7D",X"6A",X"C8",
		X"3E",X"26",X"F3",X"6F",X"5E",X"86",X"01",X"BD",X"E0",X"7D",X"FC",X"EF",X"BA",X"ED",X"C8",X"5A",
		X"A6",X"C8",X"5E",X"27",X"40",X"7A",X"B8",X"21",X"AE",X"C8",X"22",X"AE",X"88",X"14",X"A6",X"06",
		X"4A",X"26",X"32",X"86",X"01",X"BD",X"E0",X"7D",X"10",X"8E",X"64",X"74",X"86",X"00",X"5F",X"BD",
		X"E0",X"63",X"25",X"EF",X"86",X"1E",X"A7",X"28",X"8E",X"9E",X"55",X"A6",X"51",X"81",X"01",X"27",
		X"03",X"8E",X"9F",X"66",X"AF",X"29",X"AE",X"C8",X"22",X"BD",X"11",X"29",X"BD",X"3B",X"E7",X"BD",
		X"63",X"6F",X"7E",X"E0",X"69",X"0A",X"90",X"86",X"1E",X"BD",X"E0",X"7D",X"A6",X"C8",X"5E",X"27",
		X"08",X"AE",X"C8",X"22",X"BD",X"11",X"29",X"27",X"E3",X"BD",X"59",X"BF",X"7E",X"5A",X"B3",X"96",
		X"49",X"27",X"06",X"B6",X"CC",X"19",X"44",X"25",X"01",X"39",X"35",X"06",X"86",X"90",X"1F",X"31",
		X"BD",X"64",X"68",X"CC",X"03",X"84",X"ED",X"C8",X"37",X"8E",X"64",X"05",X"AF",X"C8",X"33",X"96",
		X"31",X"9A",X"40",X"27",X"73",X"B6",X"C9",X"86",X"84",X"C0",X"27",X"0D",X"F6",X"CC",X"07",X"C4",
		X"0F",X"C1",X"09",X"27",X"63",X"D6",X"E1",X"26",X"5F",X"BD",X"63",X"EE",X"AC",X"C8",X"33",X"27",
		X"18",X"34",X"12",X"AE",X"C8",X"33",X"A6",X"84",X"AE",X"01",X"5F",X"BD",X"E0",X"25",X"CC",X"03",
		X"84",X"ED",X"C8",X"37",X"35",X"12",X"AF",X"C8",X"33",X"A6",X"84",X"AE",X"01",X"10",X"AE",X"C8",
		X"22",X"E6",X"A8",X"1F",X"10",X"AE",X"C8",X"37",X"27",X"0C",X"31",X"3F",X"10",X"AF",X"C8",X"37",
		X"26",X"01",X"5F",X"BD",X"E0",X"25",X"86",X"01",X"BD",X"E0",X"7D",X"7E",X"63",X"8F",X"8E",X"64",
		X"02",X"D6",X"E1",X"26",X"0C",X"F6",X"CC",X"07",X"C4",X"0F",X"C1",X"09",X"27",X"03",X"8E",X"64",
		X"05",X"39",X"A2",X"2C",X"10",X"A1",X"2C",X"10",X"AE",X"C8",X"33",X"A6",X"84",X"AE",X"01",X"5F",
		X"BD",X"E0",X"25",X"96",X"31",X"9A",X"40",X"27",X"4C",X"8E",X"CC",X"06",X"BD",X"00",X"24",X"81",
		X"09",X"27",X"0F",X"86",X"99",X"9B",X"E1",X"19",X"97",X"E1",X"8E",X"CD",X"00",X"BD",X"00",X"2D",
		X"0C",X"6E",X"C6",X"0A",X"BD",X"00",X"1E",X"C6",X"0B",X"BD",X"00",X"1E",X"86",X"90",X"1F",X"31",
		X"BD",X"64",X"68",X"D6",X"4A",X"BD",X"00",X"48",X"96",X"4A",X"8B",X"99",X"19",X"AE",X"C8",X"22",
		X"AE",X"88",X"14",X"A7",X"05",X"E7",X"06",X"BD",X"11",X"3B",X"B6",X"B8",X"30",X"2F",X"06",X"BD",
		X"59",X"BF",X"7E",X"5A",X"B3",X"7E",X"E0",X"69",X"1F",X"89",X"E8",X"11",X"E7",X"11",X"AE",X"88",
		X"44",X"2B",X"F5",X"39",X"8E",X"00",X"70",X"6A",X"48",X"27",X"0C",X"96",X"68",X"2A",X"08",X"96",
		X"31",X"9A",X"40",X"26",X"04",X"6F",X"48",X"6F",X"4A",X"EC",X"49",X"BD",X"E0",X"56",X"86",X"02",
		X"BD",X"E0",X"7D",X"A6",X"48",X"26",X"DD",X"0A",X"90",X"7E",X"E0",X"69",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FE",X"FF",X"FE",X"FF",X"00",X"FF",X"FF",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"06",X"07",X"08",X"00",X"09",X"00",X"00",X"00",X"0A",X"00",X"00",X"02",
		X"00",X"04",X"00",X"00",X"00",X"06",X"00",X"02",X"04",X"00",X"06",X"00",X"00",X"00",X"08",X"00",
		X"00",X"FF",X"FF",X"FF",X"C0",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"0B",X"16",X"00",X"21",X"00",X"00",X"00",X"2C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FE",X"03",X"00",X"F4",X"FF",X"FF",X"FF",X"FF",X"00",X"1B",X"F9",
		X"FE",X"FD",X"F4",X"00",X"FF",X"C0",X"FF",X"00",X"00",X"1A",X"F9",X"02",X"03",X"0C",X"00",X"00",
		X"40",X"01",X"00",X"00",X"1C",X"07",X"02",X"FD",X"00",X"0C",X"00",X"01",X"00",X"01",X"00",X"1D",
		X"07",X"FD",X"01",X"FD",X"F9",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FD",X"FF",X"F9",X"FD",
		X"FF",X"C0",X"FF",X"00",X"00",X"00",X"00",X"03",X"01",X"07",X"03",X"00",X"40",X"01",X"00",X"00",
		X"00",X"00",X"03",X"FF",X"03",X"07",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FE",X"03",X"04",
		X"F8",X"FF",X"FF",X"FF",X"FF",X"02",X"00",X"00",X"FE",X"FD",X"F8",X"04",X"FF",X"C0",X"FF",X"00",
		X"02",X"00",X"00",X"02",X"03",X"08",X"FC",X"00",X"40",X"01",X"00",X"FE",X"00",X"00",X"02",X"FD",
		X"FC",X"08",X"00",X"01",X"00",X"01",X"FE",X"00",X"00",X"FD",X"03",X"01",X"F5",X"FF",X"FF",X"FF",
		X"FF",X"04",X"00",X"00",X"FD",X"FD",X"F5",X"01",X"FF",X"C0",X"FF",X"00",X"04",X"00",X"00",X"03",
		X"03",X"0B",X"FF",X"00",X"40",X"01",X"00",X"FC",X"00",X"00",X"03",X"FD",X"FF",X"0B",X"00",X"01",
		X"00",X"01",X"FC",X"00",X"00",X"B6",X"C9",X"86",X"F6",X"C9",X"85",X"C4",X"C7",X"CA",X"30",X"F7",
		X"C9",X"85",X"F6",X"C9",X"84",X"20",X"0F",X"B6",X"C9",X"86",X"44",X"F6",X"C9",X"85",X"CA",X"38",
		X"F7",X"C9",X"85",X"F6",X"C9",X"84",X"A7",X"C8",X"12",X"B6",X"C9",X"80",X"2B",X"07",X"53",X"C4",
		X"F0",X"27",X"50",X"20",X"0B",X"6F",X"C8",X"12",X"53",X"C4",X"F0",X"27",X"46",X"6C",X"C8",X"12",
		X"8E",X"66",X"27",X"A6",X"C8",X"21",X"26",X"0F",X"1F",X"98",X"A4",X"C8",X"5F",X"27",X"08",X"44",
		X"44",X"44",X"44",X"6D",X"86",X"2B",X"2A",X"A6",X"C8",X"5F",X"34",X"02",X"84",X"0F",X"A7",X"C8",
		X"5F",X"35",X"02",X"EA",X"C8",X"5F",X"E7",X"C8",X"5F",X"34",X"02",X"E8",X"E0",X"C4",X"F0",X"27",
		X"15",X"E4",X"C8",X"5F",X"26",X"03",X"E6",X"C8",X"5F",X"54",X"54",X"54",X"54",X"A6",X"85",X"2B",
		X"02",X"1F",X"89",X"E7",X"C8",X"21",X"39",X"FF",X"FF",X"FF",X"01",X"FF",X"04",X"00",X"01",X"FF",
		X"00",X"02",X"02",X"08",X"04",X"08",X"00",X"6D",X"C8",X"3B",X"27",X"03",X"6A",X"C8",X"3B",X"E6",
		X"C8",X"21",X"27",X"03",X"E7",X"C8",X"10",X"58",X"8E",X"64",X"CF",X"AE",X"85",X"AF",X"C8",X"18",
		X"43",X"A4",X"C8",X"12",X"84",X"01",X"26",X"0D",X"E6",X"C8",X"12",X"C4",X"01",X"27",X"05",X"E6",
		X"C8",X"3B",X"27",X"01",X"39",X"86",X"06",X"A7",X"C8",X"3B",X"1F",X"32",X"10",X"AE",X"A8",X"44",
		X"2A",X"07",X"A6",X"A8",X"3E",X"26",X"F5",X"20",X"16",X"1F",X"31",X"AE",X"88",X"44",X"E6",X"88",
		X"3E",X"1F",X"12",X"AE",X"88",X"44",X"2A",X"07",X"E1",X"88",X"3E",X"25",X"F6",X"20",X"EF",X"86",
		X"40",X"A7",X"A8",X"3E",X"1A",X"F0",X"CC",X"01",X"16",X"FD",X"C8",X"86",X"30",X"48",X"BF",X"C8",
		X"82",X"30",X"28",X"BF",X"C8",X"84",X"7F",X"C8",X"80",X"1C",X"EF",X"EC",X"5A",X"ED",X"3A",X"EC",
		X"5C",X"ED",X"3C",X"EC",X"5E",X"ED",X"3E",X"A6",X"42",X"A7",X"22",X"FC",X"EF",X"C0",X"ED",X"A8",
		X"5A",X"AE",X"A8",X"14",X"A6",X"89",X"91",X"02",X"44",X"44",X"84",X"3C",X"8B",X"0E",X"A7",X"A8",
		X"5E",X"A6",X"A8",X"10",X"A7",X"A8",X"21",X"8E",X"77",X"5A",X"A6",X"31",X"4A",X"27",X"03",X"8E",
		X"77",X"5D",X"BD",X"E0",X"75",X"39",X"BD",X"67",X"5A",X"86",X"01",X"BD",X"E0",X"7D",X"A6",X"5E",
		X"27",X"F7",X"6A",X"C8",X"3E",X"2F",X"5B",X"E6",X"C8",X"21",X"8E",X"64",X"E1",X"E6",X"85",X"8E",
		X"64",X"EA",X"3A",X"E6",X"02",X"EB",X"02",X"1D",X"E3",X"4C",X"ED",X"4C",X"E6",X"03",X"EB",X"03",
		X"1D",X"E3",X"4E",X"ED",X"4E",X"E6",X"08",X"EB",X"08",X"EB",X"42",X"E7",X"42",X"EC",X"84",X"AB",
		X"84",X"EB",X"01",X"AB",X"5E",X"A7",X"5E",X"1D",X"E3",X"5A",X"ED",X"5A",X"EC",X"04",X"E3",X"C8",
		X"14",X"ED",X"C8",X"14",X"EC",X"06",X"E3",X"C8",X"16",X"ED",X"C8",X"16",X"ED",X"C8",X"1C",X"ED",
		X"C8",X"1A",X"BD",X"67",X"B6",X"2A",X"0B",X"BD",X"68",X"23",X"8E",X"66",X"F2",X"86",X"01",X"7E",
		X"E0",X"6C",X"1F",X"31",X"BD",X"67",X"AD",X"7E",X"66",X"E9",X"6F",X"5E",X"6F",X"C8",X"3E",X"6F",
		X"C8",X"3B",X"BD",X"E0",X"B0",X"25",X"03",X"BD",X"E0",X"80",X"6F",X"C8",X"57",X"CC",X"00",X"00",
		X"A7",X"48",X"A7",X"C8",X"42",X"ED",X"4A",X"ED",X"C8",X"46",X"FC",X"91",X"00",X"58",X"49",X"58",
		X"49",X"34",X"02",X"FC",X"91",X"00",X"D3",X"64",X"58",X"49",X"58",X"49",X"35",X"04",X"ED",X"C8",
		X"33",X"CC",X"0C",X"0C",X"ED",X"C8",X"54",X"86",X"04",X"A7",X"C8",X"56",X"AE",X"C8",X"22",X"EC",
		X"88",X"10",X"ED",X"C8",X"2D",X"FC",X"EF",X"C0",X"ED",X"C8",X"5A",X"1F",X"31",X"6F",X"1E",X"6F",
		X"88",X"3E",X"6F",X"88",X"3B",X"39",X"EC",X"5A",X"2B",X"67",X"83",X"01",X"40",X"22",X"62",X"EC",
		X"C8",X"33",X"E1",X"C8",X"16",X"22",X"5A",X"E1",X"C8",X"17",X"22",X"55",X"A1",X"C8",X"16",X"25",
		X"50",X"A1",X"C8",X"17",X"25",X"4B",X"10",X"AE",X"C8",X"14",X"E6",X"A9",X"91",X"02",X"2F",X"3E",
		X"54",X"54",X"C4",X"3C",X"E0",X"42",X"C0",X"08",X"2E",X"37",X"E6",X"A9",X"9A",X"42",X"27",X"2E",
		X"C5",X"F0",X"26",X"16",X"E1",X"C8",X"11",X"27",X"25",X"BD",X"51",X"50",X"AE",X"84",X"2A",X"1E",
		X"A6",X"88",X"51",X"2F",X"19",X"BD",X"51",X"E9",X"20",X"14",X"BD",X"51",X"50",X"AE",X"84",X"2A",
		X"0D",X"A6",X"88",X"51",X"2F",X"08",X"BD",X"51",X"E9",X"24",X"03",X"86",X"01",X"39",X"86",X"FF",
		X"39",X"4F",X"39",X"AE",X"C8",X"2D",X"A6",X"C8",X"10",X"10",X"8E",X"68",X"36",X"E6",X"A6",X"3A",
		X"AF",X"C8",X"29",X"BD",X"E0",X"88",X"39",X"00",X"02",X"00",X"04",X"00",X"00",X"00",X"06",X"8B",
		X"0C",X"91",X"B6",X"26",X"03",X"7E",X"E0",X"A1",X"39",X"BE",X"B8",X"35",X"27",X"0E",X"A6",X"88",
		X"3E",X"2F",X"04",X"8D",X"1D",X"25",X"5C",X"AE",X"88",X"44",X"2B",X"F2",X"BE",X"B8",X"37",X"27",
		X"0E",X"A6",X"88",X"3E",X"2F",X"04",X"8D",X"0A",X"25",X"49",X"AE",X"88",X"44",X"2B",X"F2",X"1C",
		X"FE",X"39",X"EC",X"4C",X"A3",X"0C",X"2A",X"04",X"43",X"50",X"82",X"FF",X"E0",X"C8",X"54",X"82",
		X"00",X"E0",X"88",X"54",X"82",X"00",X"2A",X"29",X"EC",X"4E",X"A3",X"0E",X"2A",X"04",X"43",X"50",
		X"82",X"FF",X"E0",X"C8",X"55",X"82",X"00",X"E0",X"88",X"55",X"82",X"00",X"2A",X"13",X"E6",X"02",
		X"CB",X"04",X"E0",X"42",X"2A",X"01",X"50",X"E0",X"C8",X"56",X"C0",X"04",X"2A",X"03",X"1A",X"01",
		X"39",X"1C",X"FE",X"39",X"F6",X"C9",X"85",X"C4",X"C7",X"CA",X"30",X"20",X"05",X"F6",X"C9",X"85",
		X"CA",X"38",X"F7",X"C9",X"85",X"F6",X"C9",X"84",X"53",X"8E",X"66",X"27",X"C4",X"0F",X"27",X"3D",
		X"E4",X"C8",X"24",X"27",X"32",X"A6",X"43",X"26",X"0B",X"1F",X"98",X"A4",X"C8",X"20",X"27",X"04",
		X"6D",X"86",X"2B",X"1C",X"1F",X"98",X"E8",X"C8",X"20",X"C4",X"0F",X"27",X"1A",X"34",X"02",X"E4",
		X"E0",X"26",X"07",X"E6",X"C8",X"20",X"26",X"02",X"1F",X"89",X"C4",X"0F",X"A6",X"85",X"2B",X"02",
		X"1F",X"89",X"E4",X"C8",X"24",X"26",X"06",X"E6",X"C8",X"20",X"E4",X"C8",X"24",X"E7",X"43",X"27",
		X"03",X"E7",X"C8",X"20",X"39",X"EC",X"C8",X"16",X"58",X"58",X"44",X"56",X"44",X"56",X"B3",X"91",
		X"00",X"ED",X"C8",X"14",X"20",X"1C",X"EC",X"C8",X"16",X"58",X"58",X"44",X"56",X"44",X"56",X"B3",
		X"91",X"00",X"ED",X"C8",X"14",X"8E",X"91",X"02",X"30",X"8B",X"A6",X"84",X"84",X"E0",X"44",X"44",
		X"A7",X"42",X"A6",X"C8",X"16",X"C6",X"18",X"3D",X"ED",X"4C",X"A6",X"C8",X"17",X"C6",X"18",X"3D",
		X"C3",X"00",X"0C",X"ED",X"4E",X"A6",X"C8",X"17",X"C6",X"06",X"3D",X"34",X"06",X"A6",X"C8",X"16",
		X"C6",X"06",X"3D",X"A3",X"E1",X"C3",X"00",X"90",X"ED",X"5A",X"6F",X"5C",X"A6",X"C8",X"16",X"AB",
		X"C8",X"17",X"C6",X"04",X"3D",X"E0",X"42",X"82",X"00",X"C3",X"FF",X"9F",X"34",X"0E",X"AE",X"C8",
		X"2F",X"30",X"1E",X"86",X"05",X"BD",X"E0",X"83",X"A7",X"62",X"4F",X"E3",X"E1",X"ED",X"5D",X"6F",
		X"5F",X"35",X"04",X"1D",X"E3",X"5A",X"ED",X"5A",X"39",X"0F",X"09",X"06",X"00",X"06",X"00",X"00",
		X"00",X"09",X"34",X"32",X"B6",X"B7",X"73",X"10",X"26",X"00",X"84",X"10",X"8E",X"6A",X"3C",X"86",
		X"06",X"C6",X"FF",X"BD",X"E0",X"63",X"25",X"77",X"A6",X"42",X"A0",X"C8",X"46",X"AE",X"C8",X"14",
		X"AF",X"A8",X"14",X"E6",X"89",X"91",X"02",X"2E",X"02",X"8B",X"08",X"A7",X"A8",X"35",X"A6",X"42",
		X"80",X"04",X"A7",X"22",X"CC",X"0C",X"0C",X"ED",X"A8",X"54",X"86",X"04",X"A7",X"A8",X"56",X"CC",
		X"00",X"00",X"ED",X"2A",X"A6",X"C8",X"11",X"A7",X"A8",X"11",X"CC",X"00",X"00",X"ED",X"A8",X"31",
		X"A6",X"C8",X"21",X"A7",X"A8",X"21",X"A6",X"43",X"A7",X"23",X"EC",X"5D",X"ED",X"3D",X"EC",X"5A",
		X"ED",X"3A",X"EC",X"C8",X"16",X"ED",X"A8",X"16",X"ED",X"A8",X"1C",X"ED",X"A8",X"1A",X"EC",X"4C",
		X"ED",X"2C",X"EC",X"4E",X"ED",X"2E",X"CC",X"02",X"D4",X"ED",X"A8",X"2D",X"C3",X"00",X"02",X"ED",
		X"A8",X"29",X"8E",X"77",X"99",X"BD",X"6A",X"33",X"E6",X"A8",X"35",X"1C",X"FE",X"35",X"B2",X"1A",
		X"01",X"35",X"B2",X"96",X"B5",X"27",X"02",X"30",X"03",X"7E",X"E0",X"75",X"BD",X"E0",X"80",X"FC",
		X"EF",X"C6",X"ED",X"C8",X"5A",X"BD",X"6A",X"BB",X"BD",X"6A",X"75",X"24",X"F8",X"27",X"1E",X"86",
		X"03",X"A7",X"C8",X"21",X"8E",X"77",X"9F",X"BD",X"6A",X"33",X"AE",X"C8",X"29",X"30",X"02",X"AF",
		X"C8",X"29",X"BD",X"6A",X"BB",X"BD",X"6A",X"BB",X"6A",X"C8",X"21",X"2E",X"ED",X"6F",X"5E",X"BD",
		X"6A",X"BB",X"7E",X"E0",X"69",X"B6",X"B7",X"73",X"26",X"3C",X"AE",X"C8",X"14",X"E6",X"89",X"9A",
		X"42",X"C4",X"0F",X"27",X"11",X"BD",X"51",X"50",X"AE",X"84",X"2A",X"0A",X"A6",X"88",X"51",X"2F",
		X"05",X"BD",X"51",X"84",X"25",X"20",X"BD",X"68",X"49",X"25",X"1B",X"6C",X"5E",X"6A",X"42",X"6A",
		X"C8",X"35",X"2F",X"03",X"1C",X"FE",X"39",X"AE",X"C8",X"14",X"A6",X"89",X"91",X"02",X"84",X"0F",
		X"26",X"04",X"4F",X"1A",X"01",X"39",X"86",X"01",X"1A",X"01",X"39",X"BD",X"E0",X"88",X"86",X"01",
		X"7E",X"E0",X"7D",X"34",X"36",X"B6",X"B7",X"73",X"10",X"26",X"00",X"DC",X"10",X"8E",X"6B",X"AC",
		X"A6",X"C8",X"13",X"10",X"27",X"00",X"04",X"10",X"8E",X"6B",X"B7",X"CC",X"06",X"FF",X"BD",X"E0",
		X"78",X"10",X"25",X"00",X"C3",X"0C",X"90",X"A6",X"42",X"8B",X"04",X"A7",X"22",X"A7",X"A8",X"35",
		X"8B",X"0E",X"A7",X"A8",X"12",X"6F",X"A8",X"3E",X"CC",X"0C",X"0C",X"ED",X"A8",X"54",X"86",X"04",
		X"A7",X"A8",X"56",X"AE",X"C8",X"14",X"E6",X"89",X"91",X"02",X"54",X"54",X"C4",X"3C",X"CB",X"0E",
		X"E7",X"A8",X"5E",X"CC",X"00",X"00",X"ED",X"2A",X"A6",X"C8",X"11",X"A7",X"A8",X"11",X"CC",X"00",
		X"00",X"ED",X"A8",X"31",X"A6",X"C8",X"21",X"A7",X"A8",X"21",X"8E",X"64",X"E1",X"E6",X"86",X"8E",
		X"64",X"EA",X"3A",X"E6",X"84",X"EB",X"84",X"1D",X"E3",X"5D",X"ED",X"3D",X"E6",X"01",X"EB",X"01",
		X"1D",X"E3",X"5A",X"ED",X"3A",X"EC",X"06",X"E3",X"C8",X"16",X"ED",X"A8",X"16",X"ED",X"A8",X"1C",
		X"ED",X"A8",X"1A",X"EC",X"04",X"E3",X"C8",X"14",X"ED",X"A8",X"14",X"E6",X"02",X"EB",X"02",X"1D",
		X"E3",X"4C",X"ED",X"2C",X"E6",X"03",X"EB",X"03",X"1D",X"E3",X"4E",X"ED",X"2E",X"CC",X"02",X"88",
		X"ED",X"A8",X"2D",X"A6",X"C8",X"13",X"A7",X"A8",X"13",X"27",X"1D",X"A6",X"43",X"8E",X"69",X"99",
		X"E6",X"86",X"E5",X"C8",X"21",X"26",X"11",X"8E",X"64",X"E1",X"E6",X"86",X"8E",X"64",X"EA",X"3A",
		X"EC",X"04",X"ED",X"A8",X"31",X"6F",X"A8",X"13",X"6F",X"C8",X"5E",X"6F",X"C8",X"48",X"8E",X"77",
		X"AE",X"BD",X"E0",X"75",X"1C",X"FE",X"35",X"B6",X"1A",X"01",X"35",X"B6",X"BD",X"E0",X"80",X"FC",
		X"EF",X"C0",X"ED",X"C8",X"5A",X"20",X"2F",X"BD",X"E0",X"80",X"FC",X"EF",X"C0",X"ED",X"C8",X"5A",
		X"BD",X"6C",X"1C",X"25",X"24",X"BD",X"72",X"8A",X"EC",X"04",X"E3",X"C8",X"14",X"ED",X"C8",X"14",
		X"EC",X"06",X"E3",X"C8",X"16",X"ED",X"C8",X"16",X"ED",X"C8",X"1C",X"ED",X"C8",X"1A",X"BD",X"6C",
		X"ED",X"2A",X"16",X"BD",X"6C",X"D4",X"BD",X"6C",X"1C",X"25",X"25",X"BD",X"72",X"8A",X"BD",X"6C",
		X"ED",X"2A",X"06",X"BD",X"6C",X"D4",X"7E",X"6B",X"C0",X"27",X"15",X"C1",X"02",X"22",X"11",X"8E",
		X"77",X"60",X"BD",X"E0",X"75",X"86",X"1E",X"A7",X"5F",X"BD",X"6C",X"D4",X"6A",X"5F",X"2E",X"F9",
		X"6F",X"5E",X"86",X"01",X"BD",X"E0",X"7D",X"0A",X"90",X"7E",X"E0",X"69",X"B6",X"B7",X"73",X"26",
		X"52",X"BD",X"68",X"49",X"25",X"4D",X"AE",X"C8",X"14",X"8C",X"09",X"40",X"24",X"1C",X"A6",X"89",
		X"91",X"02",X"2F",X"16",X"44",X"44",X"84",X"3C",X"A7",X"C8",X"35",X"A6",X"42",X"8B",X"08",X"2B",
		X"32",X"A1",X"C8",X"35",X"2E",X"4B",X"27",X"2E",X"2D",X"29",X"A6",X"C8",X"21",X"8E",X"64",X"E1",
		X"E6",X"86",X"8E",X"64",X"EA",X"3A",X"EC",X"04",X"E3",X"C8",X"14",X"1F",X"01",X"8C",X"09",X"40",
		X"24",X"06",X"A6",X"89",X"91",X"02",X"2E",X"CC",X"A6",X"42",X"8B",X"10",X"2B",X"05",X"A1",X"C8",
		X"35",X"2E",X"1E",X"7E",X"6C",X"D1",X"E6",X"C8",X"12",X"E0",X"C8",X"35",X"54",X"E7",X"C8",X"3E",
		X"EB",X"C8",X"35",X"E7",X"C8",X"12",X"E6",X"C8",X"3E",X"27",X"06",X"8E",X"77",X"B1",X"BD",X"E0",
		X"75",X"E6",X"C8",X"3E",X"27",X"18",X"6C",X"42",X"6C",X"C8",X"5E",X"6A",X"5E",X"6A",X"C8",X"3E",
		X"27",X"25",X"6C",X"42",X"6C",X"C8",X"5E",X"6A",X"5E",X"6A",X"C8",X"3E",X"20",X"19",X"A1",X"C8",
		X"35",X"27",X"14",X"4A",X"6A",X"42",X"6A",X"C8",X"5E",X"6C",X"5E",X"A1",X"C8",X"35",X"27",X"07",
		X"6A",X"42",X"6A",X"C8",X"5E",X"6C",X"5E",X"EC",X"5A",X"83",X"01",X"20",X"24",X"03",X"1C",X"FE",
		X"39",X"1A",X"01",X"39",X"AE",X"C8",X"2D",X"6C",X"C8",X"1E",X"A6",X"C8",X"1E",X"46",X"24",X"02",
		X"30",X"02",X"AF",X"C8",X"29",X"BD",X"E0",X"88",X"86",X"01",X"7E",X"E0",X"7D",X"10",X"AE",X"C8",
		X"14",X"10",X"8C",X"09",X"40",X"24",X"1A",X"E6",X"A9",X"91",X"02",X"2F",X"14",X"E6",X"A9",X"9A",
		X"42",X"27",X"0E",X"E1",X"C8",X"11",X"27",X"09",X"34",X"04",X"BD",X"51",X"84",X"35",X"04",X"25",
		X"2A",X"EC",X"C8",X"31",X"27",X"3C",X"E3",X"C8",X"14",X"1F",X"02",X"10",X"8C",X"09",X"40",X"24",
		X"31",X"E6",X"A9",X"91",X"02",X"2F",X"2B",X"E6",X"A9",X"9A",X"42",X"27",X"25",X"E1",X"C8",X"11",
		X"27",X"20",X"34",X"04",X"BD",X"51",X"84",X"35",X"04",X"24",X"17",X"A6",X"11",X"81",X"03",X"25",
		X"0E",X"22",X"0A",X"F6",X"B7",X"48",X"26",X"0A",X"A6",X"88",X"51",X"2F",X"05",X"4F",X"39",X"86",
		X"01",X"39",X"86",X"FF",X"39",X"B6",X"B7",X"73",X"26",X"F3",X"10",X"AE",X"C8",X"14",X"10",X"8C",
		X"09",X"40",X"24",X"24",X"E6",X"A9",X"91",X"02",X"2F",X"1E",X"54",X"54",X"C4",X"3C",X"E0",X"42",
		X"C0",X"08",X"2E",X"D9",X"E6",X"A9",X"9A",X"42",X"27",X"0E",X"E1",X"C8",X"11",X"27",X"09",X"34",
		X"04",X"BD",X"51",X"84",X"35",X"04",X"25",X"B3",X"EC",X"C8",X"31",X"27",X"C5",X"E3",X"C8",X"14",
		X"1F",X"02",X"10",X"8C",X"09",X"40",X"24",X"BA",X"E6",X"A9",X"91",X"02",X"2F",X"B4",X"54",X"54",
		X"C4",X"3C",X"E0",X"42",X"C0",X"08",X"2E",X"A5",X"7E",X"6D",X"27",X"BD",X"E0",X"80",X"FC",X"EF",
		X"C0",X"ED",X"C8",X"5A",X"20",X"34",X"BD",X"E0",X"80",X"FC",X"EF",X"C0",X"ED",X"C8",X"5A",X"6A",
		X"C8",X"12",X"2F",X"29",X"BD",X"72",X"8A",X"EC",X"04",X"E3",X"C8",X"14",X"ED",X"C8",X"14",X"EC",
		X"06",X"E3",X"C8",X"16",X"ED",X"C8",X"16",X"ED",X"C8",X"1C",X"ED",X"C8",X"1A",X"BD",X"68",X"49",
		X"25",X"33",X"BD",X"6D",X"55",X"2A",X"1B",X"BD",X"6E",X"21",X"6A",X"C8",X"12",X"2F",X"26",X"BD",
		X"72",X"8A",X"BD",X"68",X"49",X"25",X"1E",X"BD",X"6D",X"55",X"2A",X"06",X"BD",X"6E",X"21",X"7E",
		X"6D",X"BF",X"27",X"11",X"C1",X"02",X"22",X"0D",X"86",X"1E",X"A7",X"5F",X"BD",X"6E",X"21",X"6A",
		X"5F",X"2E",X"F9",X"20",X"00",X"6F",X"5E",X"86",X"01",X"BD",X"E0",X"7D",X"0A",X"90",X"7E",X"E0",
		X"69",X"AE",X"C8",X"2D",X"A6",X"C8",X"21",X"10",X"8E",X"6E",X"4A",X"A6",X"A6",X"30",X"86",X"6C",
		X"C8",X"1E",X"A6",X"C8",X"1E",X"81",X"03",X"25",X"04",X"4F",X"A7",X"C8",X"1E",X"48",X"30",X"86",
		X"AF",X"C8",X"29",X"BD",X"E0",X"88",X"86",X"01",X"7E",X"E0",X"7D",X"00",X"06",X"00",X"0C",X"00",
		X"00",X"00",X"12",X"F6",X"B7",X"73",X"10",X"26",X"00",X"92",X"6A",X"C8",X"39",X"2E",X"1E",X"A7",
		X"C8",X"39",X"BE",X"B7",X"16",X"27",X"05",X"A6",X"88",X"51",X"26",X"1C",X"BE",X"B7",X"18",X"27",
		X"05",X"A6",X"88",X"51",X"26",X"53",X"CC",X"00",X"00",X"ED",X"C8",X"33",X"39",X"AE",X"D8",X"37",
		X"2A",X"F4",X"A6",X"88",X"51",X"27",X"EF",X"39",X"EC",X"88",X"16",X"A0",X"C8",X"16",X"2A",X"01",
		X"40",X"E0",X"C8",X"17",X"2A",X"01",X"50",X"34",X"02",X"E1",X"E4",X"25",X"02",X"E7",X"E4",X"BE",
		X"B7",X"18",X"27",X"20",X"A6",X"88",X"51",X"27",X"1B",X"EC",X"88",X"16",X"A0",X"C8",X"16",X"2A",
		X"01",X"40",X"E0",X"C8",X"17",X"2A",X"01",X"50",X"34",X"02",X"E1",X"E0",X"22",X"02",X"1F",X"89",
		X"E1",X"E4",X"25",X"03",X"BE",X"B7",X"16",X"35",X"02",X"A6",X"02",X"A7",X"C8",X"35",X"A6",X"88",
		X"3A",X"A7",X"C8",X"36",X"EC",X"88",X"16",X"ED",X"C8",X"33",X"10",X"8E",X"B7",X"18",X"BC",X"B7",
		X"18",X"27",X"04",X"10",X"8E",X"B7",X"16",X"10",X"AF",X"C8",X"37",X"39",X"6F",X"C8",X"39",X"CC",
		X"6F",X"14",X"ED",X"C8",X"37",X"BE",X"B7",X"74",X"10",X"2A",X"FF",X"7A",X"CC",X"B7",X"74",X"ED",
		X"C8",X"37",X"A6",X"02",X"A7",X"C8",X"35",X"A6",X"88",X"3A",X"A7",X"C8",X"36",X"EC",X"88",X"16",
		X"ED",X"C8",X"33",X"39",X"00",X"00",X"A6",X"C8",X"20",X"A7",X"C8",X"21",X"39",X"B6",X"B8",X"31",
		X"81",X"0B",X"22",X"F2",X"AE",X"C8",X"22",X"EC",X"02",X"ED",X"C8",X"27",X"6E",X"D8",X"27",X"BD",
		X"70",X"07",X"CC",X"6F",X"50",X"ED",X"C8",X"27",X"F6",X"B8",X"72",X"E7",X"C8",X"12",X"BD",X"E0",
		X"72",X"48",X"B1",X"B8",X"69",X"25",X"09",X"CC",X"70",X"FC",X"ED",X"C8",X"27",X"7E",X"70",X"FC",
		X"EC",X"C8",X"33",X"27",X"09",X"6D",X"C8",X"12",X"2F",X"0A",X"6A",X"C8",X"12",X"39",X"C6",X"1E",
		X"E7",X"C8",X"12",X"39",X"BD",X"75",X"32",X"E6",X"84",X"E7",X"C8",X"21",X"81",X"07",X"22",X"ED",
		X"86",X"13",X"34",X"02",X"B6",X"B7",X"73",X"10",X"26",X"00",X"88",X"10",X"8E",X"6D",X"AB",X"A6",
		X"C8",X"13",X"27",X"04",X"10",X"8E",X"6D",X"B6",X"CC",X"06",X"FF",X"BD",X"E0",X"78",X"25",X"73",
		X"0C",X"90",X"EC",X"5A",X"ED",X"3A",X"EC",X"5D",X"ED",X"3D",X"A6",X"42",X"8B",X"04",X"A7",X"22",
		X"EC",X"C8",X"16",X"ED",X"A8",X"16",X"ED",X"A8",X"1C",X"ED",X"A8",X"1A",X"CC",X"0C",X"0C",X"ED",
		X"A8",X"54",X"86",X"04",X"A7",X"A8",X"56",X"AE",X"C8",X"14",X"AF",X"A8",X"14",X"A6",X"89",X"91",
		X"02",X"44",X"44",X"84",X"3C",X"8B",X"0E",X"A7",X"A8",X"5E",X"EC",X"4C",X"ED",X"2C",X"EC",X"4E",
		X"ED",X"2E",X"A6",X"C8",X"21",X"A7",X"A8",X"21",X"CC",X"02",X"2C",X"ED",X"A8",X"2D",X"A6",X"C8",
		X"11",X"A7",X"A8",X"11",X"A6",X"E4",X"A7",X"A8",X"12",X"8E",X"77",X"C9",X"B6",X"B7",X"48",X"27",
		X"03",X"8E",X"77",X"CC",X"BD",X"E0",X"75",X"AE",X"C8",X"22",X"EC",X"02",X"ED",X"C8",X"27",X"1C",
		X"FE",X"35",X"82",X"1A",X"01",X"35",X"82",X"A6",X"C8",X"5F",X"26",X"19",X"B6",X"B8",X"26",X"B1",
		X"B8",X"25",X"25",X"0B",X"EC",X"E1",X"A6",X"C8",X"20",X"27",X"0A",X"A7",X"C8",X"21",X"39",X"6A",
		X"C8",X"5F",X"7C",X"B8",X"26",X"39",X"BD",X"70",X"07",X"CC",X"70",X"47",X"ED",X"C8",X"27",X"F6",
		X"B8",X"75",X"E7",X"C8",X"12",X"BD",X"E0",X"72",X"48",X"B1",X"B8",X"6C",X"25",X"09",X"CC",X"70",
		X"FC",X"ED",X"C8",X"27",X"7E",X"70",X"FC",X"EC",X"C8",X"33",X"27",X"09",X"6D",X"C8",X"12",X"2F",
		X"0A",X"6A",X"C8",X"12",X"39",X"C6",X"1E",X"E7",X"C8",X"12",X"39",X"8E",X"76",X"EF",X"A0",X"C8",
		X"16",X"2A",X"04",X"40",X"30",X"88",X"10",X"E0",X"C8",X"17",X"2A",X"03",X"50",X"30",X"08",X"34",
		X"02",X"E1",X"E0",X"25",X"04",X"1E",X"89",X"30",X"04",X"C1",X"00",X"27",X"06",X"E6",X"84",X"E7",
		X"C8",X"21",X"39",X"E6",X"84",X"E7",X"C8",X"21",X"81",X"08",X"22",X"F6",X"86",X"13",X"7E",X"6F",
		X"72",X"BD",X"70",X"07",X"CC",X"70",X"B2",X"ED",X"C8",X"27",X"F6",X"B8",X"78",X"E7",X"C8",X"12",
		X"BD",X"E0",X"72",X"48",X"B1",X"B8",X"6F",X"25",X"09",X"CC",X"70",X"FC",X"ED",X"C8",X"27",X"7E",
		X"70",X"FC",X"EC",X"C8",X"33",X"27",X"09",X"6D",X"C8",X"12",X"2F",X"0A",X"6A",X"C8",X"12",X"39",
		X"C6",X"1E",X"E7",X"C8",X"12",X"39",X"8E",X"77",X"0F",X"A0",X"C8",X"16",X"2A",X"04",X"40",X"30",
		X"88",X"10",X"E0",X"C8",X"17",X"2A",X"03",X"50",X"30",X"08",X"34",X"02",X"E1",X"E0",X"25",X"04",
		X"1E",X"89",X"30",X"04",X"C1",X"00",X"27",X"06",X"E6",X"84",X"E7",X"C8",X"21",X"39",X"E6",X"84",
		X"E7",X"C8",X"21",X"81",X"08",X"22",X"F6",X"86",X"13",X"7E",X"6F",X"72",X"EC",X"C8",X"33",X"27",
		X"22",X"6D",X"C8",X"12",X"2F",X"04",X"6A",X"C8",X"12",X"39",X"BD",X"71",X"C4",X"25",X"14",X"81",
		X"09",X"22",X"F6",X"AE",X"D8",X"37",X"86",X"04",X"AB",X"02",X"A0",X"42",X"2D",X"EB",X"86",X"13",
		X"7E",X"6F",X"72",X"86",X"1E",X"A7",X"C8",X"12",X"6A",X"C8",X"3B",X"A6",X"C8",X"3B",X"40",X"85",
		X"07",X"26",X"24",X"44",X"44",X"44",X"81",X"08",X"2D",X"04",X"4F",X"6F",X"C8",X"3B",X"8E",X"71",
		X"6A",X"E6",X"C8",X"21",X"A6",X"86",X"27",X"0C",X"2A",X"05",X"8E",X"71",X"61",X"20",X"03",X"8E",
		X"71",X"58",X"E6",X"85",X"E7",X"C8",X"21",X"39",X"02",X"02",X"08",X"00",X"01",X"00",X"00",X"00",
		X"04",X"04",X"04",X"01",X"00",X"08",X"00",X"00",X"00",X"02",X"00",X"00",X"01",X"FF",X"00",X"00",
		X"FF",X"01",X"10",X"8E",X"72",X"18",X"AE",X"D8",X"37",X"2A",X"46",X"A6",X"88",X"51",X"27",X"41",
		X"EC",X"C8",X"33",X"27",X"3C",X"EC",X"88",X"16",X"A0",X"C8",X"16",X"27",X"07",X"2A",X"03",X"40",
		X"31",X"22",X"31",X"22",X"E0",X"C8",X"17",X"27",X"07",X"2A",X"03",X"50",X"31",X"26",X"31",X"26",
		X"34",X"06",X"E6",X"03",X"8E",X"72",X"0F",X"E6",X"85",X"31",X"A5",X"E6",X"21",X"27",X"07",X"E6",
		X"A4",X"E7",X"C8",X"21",X"E6",X"21",X"8E",X"72",X"72",X"3A",X"35",X"06",X"AD",X"84",X"1C",X"FE",
		X"39",X"1A",X"01",X"39",X"10",X"8E",X"72",X"18",X"AE",X"D8",X"37",X"2A",X"F4",X"A6",X"88",X"51",
		X"27",X"EF",X"EC",X"C8",X"33",X"27",X"EA",X"EC",X"88",X"16",X"A0",X"C8",X"16",X"27",X"07",X"2A",
		X"03",X"40",X"31",X"22",X"31",X"22",X"E0",X"C8",X"17",X"27",X"07",X"2A",X"03",X"50",X"31",X"26",
		X"31",X"26",X"34",X"06",X"E6",X"03",X"8E",X"72",X"0F",X"E6",X"85",X"31",X"A5",X"E6",X"A4",X"E7",
		X"C8",X"21",X"E6",X"21",X"8E",X"72",X"72",X"3A",X"35",X"06",X"AD",X"84",X"1C",X"FE",X"39",X"00",
		X"12",X"24",X"00",X"36",X"00",X"00",X"00",X"48",X"02",X"00",X"04",X"09",X"02",X"09",X"08",X"07",
		X"08",X"00",X"08",X"00",X"01",X"07",X"01",X"00",X"01",X"00",X"01",X"00",X"04",X"00",X"02",X"00",
		X"08",X"0A",X"04",X"10",X"02",X"10",X"01",X"03",X"04",X"00",X"02",X"00",X"02",X"00",X"04",X"0C",
		X"02",X"05",X"08",X"00",X"08",X"0E",X"08",X"00",X"01",X"00",X"01",X"0E",X"01",X"00",X"04",X"00",
		X"04",X"05",X"02",X"0C",X"08",X"00",X"08",X"00",X"08",X"0E",X"01",X"00",X"01",X"00",X"01",X"0E",
		X"08",X"00",X"04",X"00",X"02",X"00",X"08",X"03",X"04",X"00",X"02",X"00",X"01",X"0A",X"04",X"10",
		X"02",X"10",X"86",X"7F",X"39",X"1E",X"98",X"48",X"39",X"1E",X"98",X"39",X"1E",X"98",X"44",X"39",
		X"1E",X"98",X"58",X"34",X"04",X"A1",X"E0",X"26",X"E9",X"39",X"E6",X"C8",X"21",X"8E",X"64",X"E1",
		X"E6",X"85",X"8E",X"64",X"EA",X"3A",X"E6",X"02",X"1D",X"E3",X"4C",X"ED",X"4C",X"E6",X"03",X"1D",
		X"E3",X"4E",X"ED",X"4E",X"E6",X"08",X"EB",X"42",X"E7",X"42",X"EC",X"84",X"AB",X"5E",X"A7",X"5E",
		X"1D",X"E3",X"5A",X"ED",X"5A",X"39",X"8D",X"D5",X"EC",X"04",X"E3",X"C8",X"14",X"ED",X"C8",X"14",
		X"EC",X"06",X"E3",X"C8",X"16",X"ED",X"C8",X"16",X"E3",X"4A",X"ED",X"C8",X"1C",X"EC",X"C8",X"16",
		X"A3",X"4A",X"ED",X"C8",X"1A",X"39",X"B6",X"B8",X"31",X"27",X"08",X"6F",X"43",X"B6",X"B7",X"85",
		X"7E",X"6E",X"53",X"AE",X"C8",X"22",X"EC",X"84",X"ED",X"C8",X"25",X"6E",X"D8",X"25",X"BD",X"73",
		X"DC",X"B6",X"B7",X"7D",X"26",X"15",X"10",X"8E",X"76",X"52",X"7E",X"74",X"24",X"B6",X"B7",X"83",
		X"BD",X"6E",X"53",X"26",X"06",X"6F",X"43",X"6F",X"C8",X"20",X"39",X"FC",X"B8",X"2A",X"27",X"E6",
		X"A6",X"C8",X"20",X"A1",X"43",X"27",X"09",X"43",X"A4",X"C8",X"24",X"BD",X"75",X"57",X"20",X"27",
		X"8E",X"77",X"2F",X"E6",X"C8",X"24",X"C4",X"0F",X"E6",X"85",X"26",X"23",X"A6",X"43",X"26",X"08",
		X"A6",X"C8",X"24",X"BD",X"75",X"57",X"20",X"0F",X"A4",X"C8",X"24",X"26",X"0A",X"8E",X"77",X"3F",
		X"A6",X"43",X"A6",X"86",X"A4",X"C8",X"24",X"84",X"0F",X"A7",X"43",X"A7",X"C8",X"20",X"39",X"2A",
		X"05",X"A6",X"C8",X"24",X"20",X"F1",X"8E",X"77",X"3F",X"E6",X"43",X"A6",X"85",X"A4",X"C8",X"24",
		X"BD",X"74",X"9B",X"20",X"E2",X"BD",X"73",X"DC",X"B6",X"B7",X"7E",X"26",X"1A",X"10",X"8E",X"76",
		X"56",X"7E",X"74",X"24",X"B6",X"B7",X"84",X"BD",X"6E",X"53",X"26",X"06",X"6F",X"43",X"6F",X"C8",
		X"20",X"39",X"FC",X"B8",X"2A",X"27",X"E6",X"A6",X"C8",X"20",X"A1",X"43",X"27",X"09",X"43",X"A4",
		X"C8",X"24",X"BD",X"75",X"7F",X"20",X"27",X"8E",X"77",X"2F",X"E6",X"C8",X"24",X"C4",X"0F",X"E6",
		X"85",X"26",X"23",X"A6",X"43",X"26",X"08",X"A6",X"C8",X"24",X"BD",X"75",X"7F",X"20",X"0F",X"A4",
		X"C8",X"24",X"26",X"0A",X"8E",X"77",X"3F",X"A6",X"43",X"A6",X"86",X"A4",X"C8",X"24",X"84",X"0F",
		X"A7",X"43",X"A7",X"C8",X"20",X"39",X"2A",X"05",X"A6",X"C8",X"24",X"20",X"F1",X"8E",X"77",X"3F",
		X"E6",X"43",X"A6",X"85",X"A4",X"C8",X"24",X"BD",X"74",X"9B",X"20",X"E2",X"EC",X"E1",X"ED",X"C8",
		X"25",X"6F",X"43",X"6F",X"C8",X"20",X"FC",X"B8",X"14",X"ED",X"C8",X"33",X"58",X"58",X"44",X"56",
		X"44",X"56",X"B3",X"91",X"00",X"1F",X"01",X"E6",X"89",X"90",X"C1",X"50",X"E7",X"C8",X"36",X"96",
		X"68",X"2B",X"06",X"CC",X"74",X"09",X"ED",X"C8",X"25",X"39",X"8D",X"D0",X"10",X"8E",X"76",X"5A",
		X"20",X"12",X"B6",X"B7",X"85",X"BD",X"6E",X"53",X"26",X"06",X"6F",X"43",X"6F",X"C8",X"20",X"39",
		X"10",X"8E",X"B7",X"79",X"A6",X"C8",X"20",X"A1",X"43",X"27",X"09",X"43",X"A4",X"C8",X"24",X"BD",
		X"75",X"EF",X"20",X"27",X"8E",X"77",X"2F",X"E6",X"C8",X"24",X"C4",X"0F",X"E6",X"85",X"26",X"23",
		X"A6",X"43",X"26",X"08",X"A6",X"C8",X"24",X"BD",X"75",X"EF",X"20",X"0F",X"A4",X"C8",X"24",X"26",
		X"0A",X"8E",X"77",X"3F",X"A6",X"43",X"A6",X"86",X"A4",X"C8",X"24",X"84",X"0F",X"A7",X"43",X"A7",
		X"C8",X"20",X"39",X"2A",X"05",X"A6",X"C8",X"24",X"20",X"F1",X"8E",X"77",X"3F",X"E6",X"43",X"A6",
		X"85",X"A4",X"C8",X"24",X"BD",X"75",X"EF",X"20",X"E2",X"43",X"AA",X"C8",X"41",X"43",X"26",X"0F",
		X"A6",X"C8",X"41",X"43",X"A4",X"C8",X"24",X"26",X"06",X"6F",X"C8",X"41",X"A6",X"C8",X"24",X"BD",
		X"75",X"57",X"1F",X"89",X"EA",X"C8",X"41",X"E7",X"C8",X"41",X"39",X"AE",X"C8",X"16",X"AC",X"C8",
		X"3F",X"27",X"D6",X"AC",X"C8",X"42",X"27",X"26",X"AC",X"C8",X"45",X"27",X"43",X"AC",X"C8",X"48",
		X"27",X"5F",X"BD",X"75",X"57",X"E6",X"C8",X"3E",X"CB",X"03",X"C1",X"0C",X"25",X"01",X"5F",X"E7",
		X"C8",X"3E",X"CB",X"3F",X"31",X"C5",X"AE",X"C8",X"16",X"AF",X"A4",X"A7",X"22",X"39",X"43",X"AA",
		X"C8",X"44",X"43",X"26",X"0F",X"A6",X"C8",X"44",X"43",X"A4",X"C8",X"24",X"26",X"06",X"6F",X"C8",
		X"44",X"A6",X"C8",X"24",X"BD",X"75",X"57",X"1F",X"89",X"EA",X"C8",X"44",X"E7",X"C8",X"44",X"39",
		X"43",X"AA",X"C8",X"47",X"43",X"26",X"0F",X"A6",X"C8",X"47",X"43",X"A4",X"C8",X"24",X"26",X"06",
		X"6F",X"C8",X"47",X"A6",X"C8",X"24",X"8D",X"4F",X"1F",X"89",X"EA",X"C8",X"47",X"E7",X"C8",X"47",
		X"39",X"43",X"AA",X"C8",X"4A",X"43",X"26",X"0F",X"A6",X"C8",X"4A",X"43",X"A4",X"C8",X"24",X"26",
		X"06",X"6F",X"C8",X"4A",X"A6",X"C8",X"24",X"8D",X"2E",X"1F",X"89",X"EA",X"C8",X"4A",X"E7",X"C8",
		X"4A",X"39",X"34",X"02",X"EC",X"C8",X"33",X"8E",X"76",X"CF",X"A0",X"C8",X"16",X"2A",X"04",X"40",
		X"30",X"88",X"10",X"E0",X"C8",X"17",X"2A",X"03",X"50",X"30",X"08",X"34",X"02",X"E1",X"E4",X"25",
		X"04",X"E7",X"E4",X"30",X"04",X"35",X"86",X"85",X"0F",X"27",X"15",X"E6",X"C8",X"33",X"27",X"1D",
		X"8D",X"D0",X"E5",X"80",X"26",X"14",X"E5",X"80",X"26",X"10",X"E5",X"80",X"26",X"03",X"A6",X"84",
		X"39",X"E5",X"84",X"27",X"05",X"BD",X"E0",X"72",X"25",X"F4",X"A6",X"82",X"39",X"4F",X"39",X"85",
		X"0F",X"27",X"5B",X"34",X"02",X"EC",X"C8",X"33",X"27",X"61",X"8E",X"76",X"EF",X"A0",X"C8",X"16",
		X"2A",X"04",X"40",X"30",X"88",X"10",X"E0",X"C8",X"17",X"2A",X"03",X"50",X"30",X"08",X"34",X"02",
		X"E1",X"E4",X"25",X"18",X"E7",X"E4",X"30",X"04",X"C1",X"0A",X"25",X"22",X"48",X"34",X"04",X"A1",
		X"E0",X"23",X"1B",X"BD",X"E0",X"72",X"24",X"16",X"30",X"1C",X"20",X"12",X"81",X"0A",X"25",X"0E",
		X"58",X"34",X"04",X"A1",X"E0",X"24",X"07",X"BD",X"E0",X"72",X"24",X"02",X"30",X"04",X"35",X"06",
		X"E5",X"80",X"26",X"14",X"E5",X"80",X"26",X"10",X"E5",X"80",X"26",X"03",X"A6",X"84",X"39",X"E5",
		X"84",X"27",X"05",X"BD",X"E0",X"72",X"25",X"F4",X"A6",X"82",X"39",X"35",X"02",X"4F",X"39",X"97",
		X"A6",X"AE",X"C8",X"14",X"E6",X"89",X"90",X"C1",X"2B",X"08",X"7E",X"75",X"57",X"96",X"A6",X"7E",
		X"75",X"57",X"A6",X"C8",X"3A",X"91",X"A4",X"22",X"18",X"4A",X"D6",X"9D",X"3D",X"EB",X"C8",X"36",
		X"89",X"00",X"C3",X"A3",X"81",X"1F",X"01",X"E6",X"84",X"96",X"A6",X"BD",X"76",X"5E",X"25",X"DD",
		X"39",X"8E",X"B2",X"9A",X"A6",X"86",X"4A",X"D6",X"9D",X"3D",X"34",X"04",X"E6",X"C8",X"36",X"E6",
		X"85",X"EB",X"E0",X"89",X"00",X"C3",X"A3",X"81",X"1F",X"01",X"E6",X"84",X"1F",X"98",X"84",X"CC",
		X"C4",X"33",X"44",X"44",X"58",X"58",X"34",X"02",X"EB",X"E0",X"96",X"A6",X"BD",X"76",X"5E",X"25",
		X"AC",X"39",X"3F",X"04",X"02",X"01",X"3F",X"02",X"01",X"00",X"3F",X"02",X"00",X"00",X"34",X"02",
		X"4F",X"59",X"49",X"59",X"49",X"A6",X"A6",X"97",X"A3",X"4F",X"59",X"49",X"59",X"49",X"A6",X"A6",
		X"97",X"A2",X"4F",X"59",X"49",X"59",X"49",X"A6",X"A6",X"97",X"A1",X"4F",X"59",X"49",X"59",X"49",
		X"A6",X"A6",X"97",X"A0",X"35",X"02",X"44",X"25",X"02",X"0F",X"A0",X"44",X"25",X"02",X"0F",X"A1",
		X"44",X"25",X"02",X"0F",X"A2",X"44",X"25",X"02",X"0F",X"A3",X"D6",X"A0",X"DB",X"A1",X"DB",X"A2",
		X"DB",X"A3",X"27",X"22",X"BD",X"E0",X"72",X"49",X"3D",X"1F",X"89",X"5C",X"86",X"01",X"D0",X"A0",
		X"23",X"11",X"48",X"D0",X"A1",X"23",X"0C",X"48",X"D0",X"A2",X"23",X"07",X"48",X"D0",X"A3",X"23",
		X"02",X"20",X"03",X"1C",X"FE",X"39",X"1A",X"01",X"39",X"6F",X"43",X"6F",X"C8",X"20",X"39",X"04",
		X"08",X"01",X"02",X"08",X"04",X"02",X"01",X"04",X"01",X"08",X"02",X"01",X"04",X"02",X"08",X"02",
		X"08",X"01",X"04",X"08",X"02",X"04",X"01",X"02",X"01",X"08",X"04",X"01",X"02",X"04",X"08",X"04",
		X"08",X"01",X"02",X"08",X"04",X"02",X"01",X"04",X"01",X"08",X"02",X"01",X"04",X"02",X"08",X"02",
		X"08",X"01",X"04",X"08",X"02",X"04",X"01",X"02",X"01",X"08",X"04",X"01",X"02",X"04",X"08",X"04",
		X"08",X"01",X"02",X"08",X"04",X"02",X"01",X"04",X"01",X"08",X"02",X"01",X"04",X"02",X"08",X"02",
		X"08",X"01",X"04",X"08",X"02",X"04",X"01",X"02",X"01",X"08",X"04",X"01",X"02",X"04",X"08",X"00",
		X"FF",X"FF",X"00",X"FF",X"00",X"00",X"01",X"FF",X"00",X"00",X"01",X"00",X"01",X"01",X"02",X"FF",
		X"F7",X"FB",X"FF",X"FD",X"FF",X"FF",X"FF",X"FE",X"46",X"15",X"00",X"46",X"16",X"01",X"00",X"00",
		X"00",X"00",X"00",X"01",X"50",X"2B",X"05",X"3C",X"19",X"1E",X"28",X"0D",X"1E",X"28",X"0E",X"1E",
		X"46",X"0A",X"1E",X"46",X"1B",X"1E",X"46",X"39",X"1E",X"32",X"0C",X"03",X"00",X"00",X"03",X"33",
		X"2D",X"10",X"33",X"2E",X"10",X"33",X"37",X"10",X"1D",X"11",X"02",X"29",X"11",X"02",X"1D",X"26",
		X"3C",X"29",X"26",X"3C",X"1D",X"25",X"3C",X"29",X"25",X"3C",X"1D",X"12",X"02",X"29",X"12",X"02",
		X"1D",X"13",X"02",X"29",X"13",X"02",X"00",X"00",X"02",X"1E",X"1C",X"3C",X"2A",X"1C",X"3C",X"28",
		X"0B",X"0F",X"2B",X"0B",X"0F",X"2D",X"07",X"1E",X"25",X"14",X"05",X"00",X"00",X"05",X"27",X"24",
		X"0F",X"26",X"02",X"0F",X"3C",X"08",X"1E",X"3C",X"09",X"1E",X"26",X"1A",X"06",X"00",X"1A",X"06",
		X"27",X"27",X"1E",X"27",X"3A",X"05",X"27",X"00",X"05",X"27",X"1D",X"1E",X"27",X"10",X"1E",X"3C",
		X"1E",X"0F",X"3C",X"1F",X"0F",X"3C",X"20",X"0F",X"3C",X"21",X"0F",X"3C",X"22",X"0F",X"3C",X"23",
		X"0F",X"3C",X"0F",X"28",X"29",X"04",X"1E",X"2A",X"05",X"1E",X"2B",X"06",X"1E",X"37",X"B8",X"0F",
		X"17",X"1E",X"5A",X"18",X"3C",X"25",X"2F",X"04",X"50",X"30",X"FF",X"50",X"31",X"FF",X"50",X"3B",
		X"FF",X"50",X"3C",X"FF",X"01",X"34",X"10",X"3B",X"35",X"04",X"00",X"00",X"04",X"02",X"32",X"0F",
		X"20",X"49",X"4E",X"46",X"45",X"52",X"4E",X"4F",X"20",X"28",X"43",X"29",X"20",X"31",X"39",X"38",
		X"34",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",
		X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
