library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity inferno_graph1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of inferno_graph1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"03",X"11",X"00",X"00",X"21",X"11",
		X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"03",X"11",X"11",X"00",X"21",X"11",X"27",
		X"00",X"11",X"11",X"70",X"00",X"11",X"11",X"00",X"03",X"11",X"11",X"00",X"21",X"11",X"27",X"00",
		X"11",X"11",X"79",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"27",X"00",X"00",
		X"11",X"70",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"27",X"00",X"00",X"00",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"20",X"00",X"00",
		X"11",X"70",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"27",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"73",X"11",X"70",X"00",X"07",X"11",X"00",X"00",X"09",X"11",X"00",X"00",X"09",X"27",X"00",
		X"00",X"08",X"79",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"03",X"11",X"20",X"00",X"21",
		X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"03",X"11",X"21",X"11",X"21",X"11",
		X"73",X"11",X"11",X"11",X"07",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"21",X"11",X"27",
		X"00",X"11",X"11",X"70",X"00",X"11",X"11",X"00",X"03",X"11",X"11",X"00",X"21",X"11",X"27",X"00",
		X"11",X"11",X"79",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"27",X"00",X"00",
		X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"21",X"11",X"20",X"00",
		X"73",X"11",X"11",X"00",X"09",X"11",X"11",X"00",X"09",X"11",X"11",X"00",X"08",X"21",X"11",X"20",
		X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"03",X"11",X"11",X"11",X"21",X"11",X"21",X"11",
		X"11",X"11",X"73",X"11",X"11",X"11",X"09",X"11",X"11",X"11",X"09",X"11",X"11",X"27",X"08",X"21",
		X"11",X"79",X"00",X"73",X"11",X"00",X"00",X"07",X"11",X"00",X"00",X"09",X"27",X"00",X"00",X"09",
		X"79",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"70",X"00",X"11",X"11",X"00",X"03",X"11",X"11",X"00",X"21",X"11",X"27",X"00",
		X"11",X"11",X"79",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"03",X"11",X"27",X"00",X"21",
		X"11",X"70",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"03",X"11",X"27",X"00",X"21",X"11",
		X"70",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"03",X"11",X"11",X"00",X"21",X"11",X"27",
		X"00",X"73",X"11",X"11",X"00",X"07",X"11",X"11",X"00",X"09",X"11",X"11",X"20",X"09",X"21",X"11",
		X"11",X"08",X"73",X"11",X"11",X"00",X"09",X"11",X"11",X"00",X"09",X"11",X"11",X"20",X"08",X"21",
		X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"03",X"11",X"21",X"11",X"21",X"11",
		X"73",X"11",X"11",X"11",X"09",X"11",X"11",X"11",X"09",X"11",X"11",X"11",X"08",X"21",X"11",X"27",
		X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"03",X"11",X"11",X"11",X"21",X"11",X"21",X"11",
		X"11",X"11",X"73",X"11",X"11",X"11",X"07",X"11",X"11",X"11",X"09",X"11",X"11",X"27",X"09",X"21",
		X"11",X"11",X"08",X"73",X"11",X"11",X"00",X"09",X"11",X"11",X"00",X"09",X"21",X"11",X"20",X"08",
		X"73",X"11",X"11",X"00",X"09",X"11",X"11",X"00",X"09",X"11",X"11",X"00",X"08",X"21",X"11",X"20",
		X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"03",X"11",X"11",X"11",X"21",X"11",X"21",X"11",
		X"11",X"11",X"73",X"11",X"11",X"11",X"07",X"11",X"11",X"11",X"09",X"11",X"11",X"27",X"09",X"21",
		X"11",X"11",X"08",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"03",X"11",X"21",X"11",X"21",X"11",
		X"73",X"11",X"11",X"11",X"09",X"11",X"11",X"11",X"09",X"11",X"11",X"11",X"08",X"21",X"11",X"27",
		X"00",X"73",X"11",X"70",X"00",X"07",X"11",X"00",X"00",X"09",X"11",X"00",X"00",X"09",X"27",X"00",
		X"00",X"08",X"79",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"03",X"11",X"00",X"00",X"21",X"11",
		X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"03",X"11",X"11",X"00",X"21",X"11",X"27",
		X"00",X"31",X"11",X"13",X"00",X"77",X"11",X"11",X"00",X"90",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"00",X"31",X"11",X"00",X"00",X"77",X"11",X"00",X"00",X"90",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"90",X"00",X"00",X"20",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"03",X"11",X"00",X"00",X"21",X"11",X"20",
		X"00",X"73",X"11",X"70",X"00",X"07",X"11",X"00",X"00",X"09",X"11",X"00",X"00",X"09",X"27",X"00",
		X"00",X"08",X"79",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"73",X"11",X"70",X"00",X"07",X"11",X"00",X"00",X"09",X"11",X"00",X"20",X"09",X"27",X"00",
		X"11",X"08",X"79",X"00",X"11",X"00",X"90",X"00",X"11",X"00",X"00",X"03",X"11",X"20",X"00",X"21",
		X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"03",X"11",X"21",X"11",X"21",X"11",
		X"73",X"11",X"11",X"11",X"07",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"21",X"11",X"27",
		X"00",X"31",X"11",X"13",X"00",X"77",X"11",X"11",X"00",X"90",X"11",X"11",X"20",X"00",X"11",X"11",
		X"11",X"00",X"31",X"11",X"11",X"00",X"77",X"11",X"11",X"00",X"90",X"11",X"11",X"20",X"00",X"11",
		X"11",X"70",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"31",X"11",X"27",X"00",X"11",X"11",
		X"79",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"31",X"11",X"13",X"00",X"11",X"11",X"70",
		X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"03",X"11",X"11",X"11",X"21",X"11",X"21",X"11",
		X"11",X"11",X"73",X"11",X"11",X"11",X"09",X"11",X"11",X"11",X"09",X"11",X"11",X"27",X"08",X"21",
		X"11",X"79",X"00",X"73",X"11",X"00",X"00",X"07",X"11",X"00",X"00",X"09",X"27",X"00",X"20",X"09",
		X"79",X"00",X"11",X"08",X"00",X"00",X"11",X"00",X"00",X"03",X"11",X"00",X"00",X"21",X"11",X"20",
		X"44",X"70",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"57",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"03",X"11",X"00",X"00",X"21",X"11",
		X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"03",X"11",X"11",X"00",X"21",X"11",X"27",
		X"00",X"31",X"11",X"13",X"00",X"77",X"11",X"11",X"00",X"90",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"00",X"31",X"11",X"00",X"00",X"77",X"11",X"00",X"00",X"90",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"46",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"70",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"57",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"70",X"00",X"00",X"44",X"70",X"00",X"00",X"44",X"70",X"00",X"00",X"57",X"21",X"00",X"00",
		X"77",X"11",X"00",X"00",X"77",X"27",X"00",X"00",X"73",X"77",X"00",X"03",X"21",X"77",X"20",X"21",
		X"79",X"73",X"70",X"11",X"90",X"21",X"70",X"11",X"90",X"11",X"73",X"11",X"80",X"27",X"21",X"11",
		X"00",X"77",X"11",X"11",X"00",X"77",X"11",X"11",X"00",X"73",X"11",X"11",X"00",X"21",X"11",X"27",
		X"00",X"11",X"11",X"70",X"00",X"11",X"11",X"70",X"03",X"11",X"11",X"70",X"21",X"11",X"27",X"54",
		X"11",X"11",X"77",X"44",X"11",X"11",X"77",X"57",X"11",X"11",X"76",X"77",X"11",X"27",X"54",X"77",
		X"11",X"79",X"79",X"76",X"11",X"00",X"90",X"54",X"11",X"00",X"90",X"44",X"27",X"00",X"80",X"57",
		X"79",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"54",
		X"44",X"70",X"00",X"00",X"44",X"70",X"00",X"00",X"44",X"70",X"00",X"00",X"57",X"21",X"00",X"00",
		X"77",X"11",X"00",X"00",X"77",X"27",X"00",X"00",X"73",X"77",X"00",X"00",X"21",X"77",X"20",X"00",
		X"79",X"73",X"70",X"00",X"90",X"21",X"70",X"00",X"90",X"11",X"70",X"00",X"80",X"27",X"20",X"00",
		X"00",X"77",X"11",X"00",X"00",X"77",X"11",X"00",X"00",X"73",X"11",X"00",X"00",X"21",X"11",X"20",
		X"00",X"73",X"11",X"70",X"00",X"09",X"11",X"70",X"00",X"09",X"11",X"70",X"00",X"08",X"27",X"54",
		X"00",X"00",X"77",X"44",X"00",X"00",X"77",X"57",X"00",X"00",X"76",X"77",X"00",X"00",X"54",X"77",
		X"00",X"00",X"79",X"76",X"00",X"00",X"90",X"54",X"00",X"00",X"90",X"44",X"00",X"00",X"80",X"57",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"54",
		X"14",X"00",X"22",X"00",X"04",X"20",X"00",X"B0",X"00",X"0E",X"CB",X"2B",X"02",X"EB",X"29",X"22",
		X"00",X"AA",X"99",X"E2",X"00",X"BA",X"17",X"B3",X"00",X"23",X"11",X"00",X"0D",X"FF",X"AA",X"09",
		X"DD",X"BB",X"AA",X"B2",X"DE",X"DD",X"33",X"23",X"E0",X"DD",X"3E",X"DB",X"EB",X"DD",X"DD",X"DD",
		X"AE",X"0D",X"DD",X"FD",X"0A",X"BB",X"C0",X"DD",X"07",X"AA",X"BB",X"C0",X"6A",X"00",X"AB",X"22",
		X"60",X"00",X"A0",X"DD",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"50",X"00",X"00",
		X"00",X"00",X"22",X"00",X"00",X"42",X"B0",X"2B",X"1D",X"20",X"9B",X"22",X"00",X"0D",X"99",X"22",
		X"00",X"FC",X"19",X"BB",X"00",X"AA",X"AA",X"0A",X"00",X"AA",X"AA",X"22",X"00",X"3F",X"3B",X"00",
		X"00",X"E2",X"22",X"22",X"0E",X"DD",X"22",X"22",X"EE",X"DD",X"22",X"D2",X"EE",X"F0",X"0E",X"F0",
		X"EA",X"D0",X"0E",X"C0",X"AB",X"00",X"0E",X"10",X"0A",X"D0",X"00",X"C0",X"67",X"B0",X"0E",X"20",
		X"60",X"AA",X"0C",X"0E",X"00",X"0A",X"4D",X"0C",X"00",X"00",X"A4",X"02",X"00",X"00",X"A0",X"DD",
		X"00",X"00",X"A0",X"44",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"50",X"00",X"00",
		X"00",X"00",X"22",X"22",X"00",X"00",X"EE",X"00",X"00",X"AF",X"C3",X"22",X"00",X"AF",X"00",X"22",
		X"1C",X"AC",X"0B",X"22",X"00",X"EC",X"22",X"AA",X"00",X"CA",X"E2",X"F0",X"00",X"AA",X"2F",X"C0",
		X"00",X"AA",X"AC",X"10",X"00",X"A2",X"AC",X"10",X"00",X"22",X"AA",X"CA",X"00",X"22",X"AA",X"20",
		X"00",X"E0",X"AA",X"D0",X"00",X"20",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"60",X"AA",X"AA",X"99",
		X"60",X"2A",X"AA",X"99",X"00",X"DA",X"AA",X"99",X"00",X"D0",X"A9",X"99",X"00",X"AD",X"99",X"99",
		X"00",X"0A",X"02",X"99",X"00",X"0A",X"C2",X"99",X"00",X"00",X"DD",X"9A",X"00",X"00",X"AD",X"AA",
		X"00",X"00",X"A0",X"D0",X"00",X"00",X"A0",X"DD",X"00",X"00",X"00",X"A4",X"50",X"00",X"00",X"0A",
		X"44",X"00",X"00",X"0A",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"50",X"00",X"00",
		X"60",X"2A",X"AA",X"FF",X"00",X"DA",X"AA",X"FF",X"00",X"D0",X"AF",X"FF",X"00",X"AD",X"FF",X"FF",
		X"00",X"0A",X"0F",X"FF",X"00",X"0A",X"C2",X"FF",X"00",X"00",X"DD",X"FF",X"00",X"00",X"AD",X"FA",
		X"00",X"00",X"A0",X"D0",X"00",X"00",X"A0",X"DD",X"00",X"00",X"00",X"A4",X"50",X"00",X"00",X"0A",
		X"44",X"00",X"00",X"0A",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"50",X"00",X"00",
		X"60",X"2A",X"AA",X"FF",X"00",X"DA",X"AA",X"EF",X"00",X"D0",X"AF",X"FF",X"00",X"AD",X"FF",X"FF",
		X"00",X"0A",X"FF",X"FF",X"00",X"0A",X"F3",X"FF",X"00",X"0F",X"FF",X"FF",X"00",X"FF",X"FF",X"FA",
		X"00",X"FF",X"FF",X"D0",X"00",X"EF",X"F3",X"DD",X"0F",X"EF",X"FF",X"A4",X"FF",X"FF",X"F0",X"0A",
		X"44",X"BF",X"00",X"0A",X"44",X"FF",X"00",X"00",X"44",X"FF",X"00",X"00",X"44",X"F0",X"00",X"00",
		X"14",X"00",X"22",X"00",X"04",X"20",X"00",X"B0",X"00",X"0E",X"22",X"2B",X"02",X"EA",X"22",X"22",
		X"00",X"AA",X"32",X"E2",X"00",X"BA",X"20",X"B3",X"00",X"23",X"D2",X"00",X"0D",X"FF",X"AA",X"09",
		X"DD",X"BB",X"AA",X"B2",X"DE",X"DD",X"33",X"23",X"E0",X"DD",X"3E",X"DB",X"EB",X"DD",X"DD",X"DD",
		X"AE",X"0D",X"DD",X"FD",X"0A",X"BB",X"C0",X"DD",X"07",X"AA",X"BB",X"C0",X"6A",X"00",X"AB",X"22",
		X"14",X"00",X"22",X"00",X"04",X"20",X"00",X"B0",X"00",X"0E",X"1B",X"2B",X"02",X"EB",X"91",X"22",
		X"00",X"AC",X"99",X"E2",X"00",X"BA",X"C9",X"B3",X"00",X"23",X"01",X"00",X"0D",X"FF",X"AA",X"09",
		X"DD",X"BB",X"AA",X"B2",X"DE",X"DD",X"33",X"23",X"E0",X"DD",X"3E",X"DB",X"EB",X"DD",X"DD",X"DD",
		X"AE",X"0D",X"DD",X"FD",X"0A",X"BB",X"C0",X"DD",X"07",X"AA",X"BB",X"C0",X"6A",X"00",X"AB",X"22",
		X"10",X"00",X"22",X"20",X"20",X"B2",X"BB",X"44",X"E0",X"22",X"CC",X"42",X"3B",X"2B",X"11",X"04",
		X"3B",X"B0",X"11",X"A0",X"E3",X"0C",X"11",X"2F",X"EE",X"00",X"CA",X"FF",X"EE",X"0A",X"AA",X"BB",
		X"FE",X"BA",X"AA",X"DD",X"DD",X"2F",X"33",X"DD",X"DD",X"EE",X"AA",X"DD",X"DD",X"BB",X"DD",X"EC",
		X"DD",X"DD",X"DD",X"0D",X"02",X"DD",X"00",X"BB",X"00",X"10",X"BB",X"A0",X"0D",X"2D",X"A0",X"A0",
		X"00",X"00",X"77",X"77",X"00",X"00",X"FF",X"F8",X"00",X"00",X"FF",X"F8",X"00",X"00",X"FF",X"F8",
		X"00",X"00",X"FF",X"F8",X"00",X"00",X"FF",X"F8",X"00",X"00",X"FF",X"F8",X"00",X"00",X"FF",X"F8",
		X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"DF",X"DF",X"00",X"00",X"DF",X"FF",
		X"00",X"00",X"DF",X"FF",X"00",X"00",X"DF",X"FF",X"00",X"00",X"DD",X"DF",X"00",X"00",X"77",X"77",
		X"77",X"77",X"77",X"77",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"DD",X"FF",X"FF",X"DD",X"DF",X"FF",X"FF",X"DF",
		X"DD",X"FF",X"FF",X"DD",X"DF",X"FF",X"FF",X"FF",X"DD",X"FF",X"FF",X"DD",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"88",X"88",X"88",X"FF",X"88",X"88",X"88",X"FF",X"88",X"88",X"88",X"FF",
		X"88",X"88",X"88",X"FF",X"88",X"88",X"88",X"FF",X"88",X"88",X"88",X"FF",X"88",X"88",X"88",X"FF",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"DF",X"DF",X"FF",X"FF",X"DF",X"DF",X"FF",X"FF",
		X"DF",X"DF",X"FF",X"FF",X"DF",X"DF",X"FF",X"FF",X"DF",X"DD",X"FF",X"FF",X"77",X"77",X"77",X"77",
		X"07",X"77",X"77",X"77",X"07",X"FF",X"88",X"88",X"07",X"FF",X"88",X"88",X"07",X"FF",X"88",X"88",
		X"07",X"FF",X"88",X"88",X"07",X"FF",X"88",X"88",X"07",X"FF",X"88",X"88",X"07",X"FF",X"88",X"88",
		X"07",X"77",X"77",X"77",X"07",X"77",X"77",X"77",X"07",X"DD",X"DF",X"FF",X"07",X"FD",X"FF",X"FF",
		X"07",X"FD",X"DF",X"FF",X"07",X"FD",X"FF",X"FF",X"07",X"DD",X"FF",X"FF",X"07",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"FF",X"FF",X"DD",X"DF",X"FF",X"FF",X"DF",X"DF",
		X"FF",X"FF",X"DF",X"DF",X"FF",X"FF",X"DF",X"DF",X"FF",X"FF",X"DD",X"DF",X"77",X"77",X"77",X"77",
		X"77",X"77",X"70",X"00",X"88",X"FF",X"70",X"00",X"88",X"FF",X"70",X"00",X"88",X"FF",X"70",X"00",
		X"88",X"FF",X"70",X"00",X"88",X"FF",X"70",X"00",X"88",X"FF",X"70",X"00",X"88",X"FF",X"70",X"00",
		X"77",X"77",X"70",X"00",X"77",X"77",X"70",X"00",X"FF",X"FF",X"70",X"00",X"FF",X"FF",X"70",X"00",
		X"FF",X"FF",X"70",X"00",X"FF",X"FF",X"70",X"00",X"FF",X"FF",X"70",X"00",X"77",X"77",X"70",X"00",
		X"44",X"70",X"00",X"64",X"44",X"00",X"00",X"77",X"44",X"00",X"00",X"90",X"57",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"03",X"11",X"00",X"00",X"21",X"11",X"20",
		X"44",X"70",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"57",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"46",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"70",X"00",X"64",X"44",X"00",X"00",X"77",X"44",X"00",X"00",X"90",X"57",X"00",X"40",X"00",
		X"79",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"06",X"44",X"00",X"00",X"54",X"44",X"50",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"06",X"44",X"44",X"44",X"54",X"44",X"54",X"44",
		X"44",X"44",X"76",X"44",X"44",X"44",X"09",X"44",X"44",X"44",X"09",X"44",X"44",X"57",X"08",X"54",
		X"44",X"44",X"00",X"64",X"44",X"44",X"00",X"77",X"44",X"44",X"00",X"90",X"54",X"44",X"50",X"00",
		X"76",X"44",X"44",X"00",X"07",X"44",X"44",X"00",X"09",X"44",X"44",X"00",X"09",X"54",X"44",X"50",
		X"08",X"44",X"44",X"70",X"00",X"44",X"44",X"00",X"06",X"44",X"44",X"00",X"54",X"44",X"57",X"00",
		X"44",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"00",X"06",X"44",X"57",X"00",X"54",
		X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"06",X"44",X"54",X"44",X"54",X"44",
		X"76",X"44",X"44",X"44",X"07",X"44",X"44",X"44",X"09",X"44",X"44",X"44",X"09",X"54",X"44",X"57",
		X"08",X"76",X"44",X"79",X"00",X"09",X"44",X"00",X"00",X"09",X"44",X"00",X"00",X"08",X"57",X"00",
		X"46",X"00",X"07",X"00",X"44",X"00",X"09",X"00",X"44",X"00",X"00",X"06",X"44",X"00",X"00",X"54",
		X"44",X"70",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"57",X"00",X"40",X"00",
		X"79",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"06",X"44",X"00",X"00",X"54",X"44",X"50",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"06",X"44",X"44",X"44",X"54",X"44",X"54",X"44",
		X"44",X"44",X"76",X"44",X"44",X"44",X"09",X"44",X"44",X"44",X"09",X"44",X"44",X"57",X"08",X"54",
		X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"54",X"44",X"50",X"00",
		X"76",X"44",X"44",X"00",X"07",X"44",X"44",X"00",X"09",X"44",X"44",X"00",X"09",X"54",X"44",X"50",
		X"08",X"44",X"44",X"70",X"00",X"44",X"44",X"00",X"06",X"44",X"44",X"00",X"54",X"44",X"57",X"00",
		X"44",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"00",X"06",X"44",X"57",X"00",X"54",
		X"44",X"44",X"00",X"64",X"44",X"44",X"00",X"77",X"44",X"44",X"00",X"90",X"54",X"44",X"50",X"00",
		X"76",X"44",X"44",X"00",X"07",X"44",X"44",X"00",X"09",X"44",X"44",X"00",X"09",X"54",X"44",X"50",
		X"08",X"44",X"44",X"70",X"00",X"44",X"44",X"00",X"06",X"44",X"44",X"00",X"54",X"44",X"57",X"00",
		X"44",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"00",X"00",X"44",X"57",X"00",X"00",
		X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"06",X"44",X"54",X"44",X"54",X"44",
		X"76",X"44",X"44",X"44",X"07",X"44",X"44",X"44",X"09",X"44",X"44",X"44",X"09",X"54",X"44",X"57",
		X"08",X"76",X"44",X"79",X"00",X"09",X"44",X"00",X"00",X"09",X"44",X"00",X"00",X"08",X"57",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"54",
		X"44",X"70",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"57",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"46",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"06",X"44",X"00",X"00",X"54",
		X"44",X"70",X"00",X"64",X"44",X"00",X"00",X"77",X"44",X"00",X"00",X"90",X"57",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"46",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"70",X"00",X"64",X"44",X"00",X"00",X"77",X"44",X"00",X"00",X"90",X"57",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"46",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"06",X"44",X"00",X"00",X"54",
		X"44",X"70",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"57",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"46",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"46",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"46",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"06",X"44",X"00",X"00",X"54",
		X"44",X"70",X"00",X"64",X"44",X"00",X"00",X"77",X"44",X"00",X"00",X"90",X"57",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"70",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"06",X"44",X"57",X"00",X"54",X"44",
		X"79",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"06",X"44",X"44",X"00",X"54",X"44",X"57",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"06",X"44",X"44",X"44",X"54",X"44",X"54",X"44",
		X"44",X"44",X"76",X"44",X"44",X"44",X"09",X"44",X"44",X"44",X"09",X"44",X"44",X"57",X"08",X"54",
		X"44",X"46",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"64",X"44",X"44",X"44",X"44",X"44",
		X"64",X"44",X"44",X"44",X"77",X"44",X"44",X"44",X"00",X"44",X"44",X"46",X"00",X"44",X"44",X"70",
		X"00",X"64",X"44",X"46",X"00",X"77",X"44",X"44",X"00",X"90",X"44",X"44",X"00",X"00",X"44",X"44",
		X"46",X"00",X"64",X"44",X"44",X"00",X"77",X"44",X"44",X"00",X"90",X"44",X"44",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"06",X"44",X"00",X"00",X"54",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"06",X"44",X"44",X"00",X"54",X"44",X"57",
		X"00",X"44",X"44",X"79",X"00",X"44",X"44",X"00",X"06",X"44",X"44",X"00",X"54",X"44",X"57",X"00",
		X"44",X"44",X"79",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"06",X"44",X"57",X"00",X"54",
		X"44",X"70",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"06",X"44",X"57",X"00",X"54",X"44",
		X"79",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"06",X"44",X"44",X"00",X"54",X"44",X"57",
		X"00",X"44",X"44",X"79",X"00",X"44",X"44",X"00",X"06",X"44",X"44",X"00",X"54",X"44",X"57",X"00",
		X"44",X"44",X"79",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"57",X"00",X"00",
		X"44",X"70",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"06",X"44",X"57",X"00",X"54",X"44",
		X"79",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"06",X"44",X"44",X"00",X"54",X"44",X"57",
		X"00",X"44",X"44",X"79",X"00",X"44",X"44",X"00",X"06",X"44",X"44",X"00",X"54",X"44",X"57",X"00",
		X"44",X"44",X"79",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"06",X"44",X"57",X"00",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"06",X"44",X"00",X"00",X"54",X"44",X"50",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"06",X"44",X"44",X"44",X"54",X"44",X"54",X"44",
		X"44",X"44",X"76",X"44",X"44",X"44",X"09",X"44",X"44",X"44",X"09",X"44",X"44",X"57",X"08",X"54",
		X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"54",X"44",X"50",X"00",
		X"76",X"44",X"44",X"00",X"07",X"44",X"44",X"00",X"09",X"44",X"44",X"00",X"09",X"54",X"44",X"50",
		X"08",X"44",X"44",X"70",X"00",X"44",X"44",X"00",X"06",X"44",X"44",X"00",X"54",X"44",X"57",X"00",
		X"44",X"44",X"77",X"00",X"44",X"44",X"09",X"00",X"44",X"44",X"00",X"00",X"44",X"57",X"00",X"00",
		X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"06",X"44",X"54",X"44",X"54",X"44",
		X"76",X"44",X"44",X"44",X"07",X"44",X"44",X"44",X"09",X"44",X"44",X"44",X"09",X"54",X"44",X"57",
		X"08",X"76",X"44",X"79",X"00",X"09",X"44",X"00",X"00",X"09",X"44",X"00",X"00",X"08",X"57",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"06",X"44",X"00",X"00",X"54",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"06",X"44",X"44",X"00",X"54",X"44",X"57",
		X"00",X"44",X"44",X"79",X"00",X"44",X"44",X"00",X"06",X"44",X"44",X"00",X"54",X"44",X"57",X"00",
		X"44",X"44",X"79",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"57",X"00",X"00",
		X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"06",X"44",X"54",X"44",X"54",X"44",
		X"76",X"44",X"44",X"44",X"09",X"44",X"44",X"44",X"09",X"44",X"44",X"44",X"08",X"54",X"44",X"57",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"06",X"44",X"44",X"44",X"54",X"44",X"54",X"44",
		X"44",X"44",X"76",X"44",X"44",X"44",X"09",X"44",X"44",X"44",X"09",X"44",X"44",X"57",X"08",X"54",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"06",X"44",X"00",X"00",X"54",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"06",X"44",X"44",X"00",X"54",X"44",X"57",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"06",X"44",X"44",X"44",X"54",X"44",X"54",X"44",
		X"44",X"44",X"76",X"44",X"44",X"44",X"09",X"44",X"44",X"44",X"09",X"44",X"44",X"57",X"08",X"54",
		X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"06",X"44",X"54",X"44",X"54",X"44",
		X"76",X"44",X"44",X"44",X"07",X"44",X"44",X"44",X"09",X"44",X"44",X"44",X"09",X"54",X"44",X"57",
		X"08",X"44",X"44",X"79",X"00",X"44",X"44",X"00",X"06",X"44",X"44",X"00",X"54",X"44",X"57",X"00",
		X"44",X"44",X"79",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"57",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"54",
		X"44",X"70",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"57",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"46",X"00",X"00",X"00",X"44",X"00",X"00",X"64",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"64",X"44",X"00",X"00",X"97",X"44",X"00",X"00",X"90",X"44",X"00",X"00",X"80",X"44",
		X"00",X"00",X"00",X"CF",X"00",X"00",X"00",X"DF",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"DF",
		X"00",X"00",X"00",X"DA",X"00",X"00",X"00",X"DA",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"D0",
		X"00",X"00",X"00",X"DB",X"00",X"00",X"00",X"D0",X"00",X"00",X"64",X"C0",X"00",X"00",X"40",X"DD",
		X"00",X"00",X"64",X"00",X"00",X"00",X"97",X"04",X"00",X"00",X"90",X"44",X"00",X"00",X"80",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"D0",X"A0",
		X"00",X"00",X"DA",X"F0",X"00",X"00",X"ED",X"EB",X"00",X"00",X"FC",X"FF",X"00",X"00",X"FE",X"DF",
		X"00",X"00",X"FD",X"CF",X"00",X"00",X"FD",X"CF",X"00",X"00",X"EB",X"FF",X"00",X"00",X"FB",X"DF",
		X"00",X"00",X"FF",X"DD",X"00",X"00",X"0F",X"FC",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"13",X"00",X"00",X"00",X"11",X"00",X"00",X"31",X"11",X"00",X"00",X"11",X"11",X"00",X"00",
		X"31",X"11",X"13",X"00",X"77",X"11",X"11",X"00",X"90",X"11",X"11",X"00",X"00",X"11",X"11",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"AD",X"00",X"00",
		X"00",X"AD",X"00",X"00",X"00",X"AD",X"00",X"00",X"00",X"AC",X"00",X"00",X"00",X"0D",X"00",X"00",
		X"00",X"AD",X"00",X"00",X"00",X"AD",X"00",X"00",X"31",X"BC",X"00",X"00",X"11",X"BD",X"00",X"00",
		X"31",X"D0",X"13",X"00",X"77",X"00",X"11",X"00",X"90",X"11",X"11",X"00",X"00",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"F0",X"00",X"00",X"EB",X"F0",X"00",X"00",X"BD",X"FA",X"00",X"00",
		X"BD",X"FF",X"00",X"00",X"FE",X"FE",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"CD",X"00",X"00",
		X"FF",X"CC",X"00",X"00",X"FF",X"EC",X"00",X"00",X"BE",X"FF",X"00",X"00",X"0F",X"FD",X"00",X"00",
		X"0F",X"DD",X"00",X"00",X"00",X"CF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"B0",
		X"00",X"00",X"00",X"3D",X"00",X"00",X"0D",X"2C",X"00",X"00",X"0D",X"33",X"00",X"00",X"00",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"00",X"DB",X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"20",X"00",X"00",X"0D",X"20",
		X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"CD",X"00",X"00",X"00",X"CD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",
		X"00",X"00",X"00",X"2D",X"00",X"00",X"00",X"CD",X"00",X"00",X"00",X"CD",X"00",X"00",X"00",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D6",X"00",X"00",X"00",X"BD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"3D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"3C",X"00",X"00",X"00",X"23",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"20",X"00",X"00",X"0D",X"33",X"00",X"00",X"02",X"C2",
		X"00",X"00",X"00",X"DC",X"00",X"00",X"00",X"DC",X"00",X"00",X"06",X"2D",X"00",X"0D",X"5F",X"FF",
		X"00",X"03",X"FD",X"FF",X"00",X"02",X"FD",X"FF",X"00",X"03",X"D3",X"FF",X"D0",X"5D",X"DF",X"57",
		X"D0",X"FD",X"FF",X"44",X"00",X"DD",X"FF",X"44",X"06",X"DD",X"FF",X"44",X"5F",X"CF",X"54",X"44",
		X"FF",X"FF",X"76",X"44",X"FF",X"FF",X"09",X"44",X"DD",X"FF",X"09",X"44",X"CF",X"57",X"08",X"54",
		X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"2D",X"00",X"03",X"0D",X"2B",X"00",X"03",X"5D",X"FF",
		X"D0",X"03",X"F3",X"FF",X"D0",X"03",X"F3",X"FF",X"00",X"0B",X"CF",X"FF",X"00",X"5D",X"DF",X"57",
		X"00",X"FD",X"FF",X"44",X"00",X"D3",X"FF",X"44",X"06",X"D3",X"FF",X"44",X"5F",X"DF",X"54",X"44",
		X"DF",X"FF",X"76",X"44",X"DD",X"FF",X"09",X"44",X"CD",X"FF",X"09",X"44",X"3F",X"57",X"08",X"54",
		X"00",X"00",X"00",X"2D",X"D0",X"00",X"0D",X"2C",X"D0",X"0D",X"0D",X"D2",X"00",X"0C",X"53",X"FF",
		X"00",X"03",X"F2",X"FF",X"00",X"0D",X"D3",X"FF",X"00",X"0D",X"CF",X"FF",X"00",X"5F",X"DF",X"57",
		X"00",X"FD",X"FF",X"44",X"00",X"DD",X"FF",X"44",X"D6",X"DF",X"FF",X"44",X"DF",X"DF",X"54",X"44",
		X"DD",X"FF",X"76",X"44",X"BD",X"FF",X"09",X"44",X"2C",X"FF",X"09",X"44",X"3F",X"57",X"08",X"54",
		X"00",X"00",X"0D",X"32",X"00",X"00",X"03",X"D2",X"00",X"00",X"02",X"D3",X"00",X"00",X"53",X"FF",
		X"00",X"00",X"FD",X"FF",X"00",X"00",X"DD",X"FF",X"00",X"06",X"CD",X"FF",X"D0",X"5F",X"DF",X"57",
		X"D0",X"FD",X"FF",X"44",X"D0",X"DD",X"FF",X"44",X"D6",X"DF",X"FF",X"44",X"BF",X"DF",X"54",X"44",
		X"2D",X"FF",X"76",X"44",X"3D",X"FF",X"09",X"44",X"2D",X"FF",X"09",X"44",X"CF",X"57",X"08",X"54",
		X"00",X"00",X"03",X"D3",X"00",X"00",X"00",X"DB",X"00",X"00",X"06",X"DD",X"00",X"00",X"5D",X"FF",
		X"00",X"00",X"FD",X"FF",X"00",X"00",X"DD",X"FF",X"00",X"06",X"CD",X"FF",X"D0",X"5D",X"DF",X"57",
		X"D0",X"FD",X"FF",X"44",X"00",X"DD",X"FF",X"44",X"26",X"DF",X"FF",X"44",X"3F",X"DF",X"54",X"44",
		X"BD",X"FF",X"76",X"44",X"DD",X"FF",X"09",X"44",X"DD",X"FF",X"09",X"44",X"DF",X"57",X"08",X"54",
		X"00",X"00",X"00",X"DC",X"00",X"00",X"00",X"DC",X"00",X"00",X"06",X"2D",X"00",X"0D",X"5F",X"FF",
		X"00",X"03",X"FD",X"FF",X"00",X"02",X"FD",X"FF",X"00",X"03",X"D3",X"FF",X"D0",X"5D",X"DF",X"57",
		X"D0",X"FD",X"FF",X"FF",X"00",X"DD",X"FF",X"FF",X"06",X"DD",X"FF",X"FF",X"5F",X"CF",X"5F",X"FF",
		X"FF",X"FF",X"76",X"FF",X"FF",X"FF",X"09",X"FF",X"DD",X"FF",X"09",X"FF",X"CF",X"57",X"08",X"5F",
		X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"2D",X"00",X"03",X"0D",X"2B",X"00",X"03",X"5D",X"FF",
		X"D0",X"03",X"F3",X"FF",X"D0",X"03",X"F3",X"FF",X"00",X"0B",X"CF",X"FF",X"00",X"5D",X"DF",X"57",
		X"00",X"FD",X"FF",X"FF",X"00",X"D3",X"FF",X"FF",X"06",X"D3",X"FF",X"FF",X"5F",X"DF",X"5F",X"FF",
		X"DF",X"FF",X"76",X"FF",X"DD",X"FF",X"09",X"FF",X"CD",X"FF",X"09",X"FF",X"3F",X"57",X"08",X"5F",
		X"00",X"00",X"00",X"2D",X"D0",X"00",X"0D",X"2C",X"D0",X"0D",X"0D",X"D2",X"00",X"0C",X"53",X"FF",
		X"00",X"03",X"F2",X"FF",X"00",X"0D",X"D3",X"FF",X"00",X"0D",X"CF",X"FF",X"00",X"5F",X"DF",X"57",
		X"00",X"FD",X"FF",X"FF",X"00",X"DD",X"FF",X"FF",X"D6",X"DF",X"FF",X"FF",X"DF",X"DF",X"5F",X"FF",
		X"DD",X"FF",X"76",X"FF",X"BD",X"FF",X"09",X"FF",X"2C",X"FF",X"09",X"FF",X"3F",X"57",X"08",X"5F",
		X"00",X"00",X"0D",X"32",X"00",X"00",X"03",X"D2",X"00",X"00",X"02",X"D3",X"00",X"00",X"53",X"FF",
		X"00",X"00",X"FD",X"FF",X"00",X"00",X"DD",X"FF",X"00",X"06",X"CD",X"FF",X"D0",X"5F",X"DF",X"57",
		X"D0",X"FD",X"FF",X"FF",X"D0",X"DD",X"FF",X"FF",X"D6",X"DF",X"FF",X"FF",X"BF",X"DF",X"5F",X"FF",
		X"2D",X"FF",X"76",X"FF",X"3D",X"FF",X"09",X"FF",X"2D",X"FF",X"09",X"FF",X"CF",X"57",X"08",X"5F",
		X"00",X"00",X"03",X"D3",X"00",X"00",X"00",X"DB",X"00",X"00",X"06",X"DD",X"00",X"00",X"5D",X"FF",
		X"00",X"00",X"FD",X"FF",X"00",X"00",X"DD",X"FF",X"00",X"06",X"CD",X"FF",X"D0",X"5D",X"DF",X"57",
		X"D0",X"FD",X"FF",X"FF",X"00",X"DD",X"FF",X"FF",X"26",X"DF",X"FF",X"FF",X"3F",X"DF",X"5F",X"FF",
		X"BD",X"FF",X"76",X"FF",X"DD",X"FF",X"09",X"FF",X"DD",X"FF",X"09",X"FF",X"DF",X"57",X"08",X"5F",
		X"00",X"00",X"00",X"DC",X"00",X"00",X"00",X"DC",X"00",X"00",X"06",X"2D",X"00",X"0D",X"5F",X"FF",
		X"00",X"03",X"FD",X"DF",X"00",X"02",X"FD",X"FF",X"00",X"03",X"D3",X"FF",X"D0",X"5D",X"DF",X"57",
		X"D0",X"FD",X"FF",X"DF",X"00",X"DD",X"FF",X"DF",X"06",X"DD",X"FF",X"DF",X"5F",X"CF",X"5F",X"BF",
		X"FF",X"FF",X"76",X"3D",X"FF",X"FF",X"0D",X"2C",X"DD",X"FF",X"0D",X"33",X"CF",X"57",X"08",X"C3",
		X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"2D",X"00",X"03",X"0D",X"2B",X"00",X"03",X"5D",X"FF",
		X"D0",X"03",X"F3",X"FF",X"D0",X"03",X"F3",X"FF",X"00",X"0B",X"CF",X"FF",X"00",X"5D",X"DF",X"5D",
		X"00",X"FD",X"FF",X"DB",X"00",X"D3",X"FF",X"BD",X"06",X"D3",X"FF",X"2F",X"5F",X"DF",X"5D",X"2F",
		X"DF",X"FF",X"76",X"CF",X"DD",X"FF",X"09",X"DD",X"CD",X"FF",X"09",X"CD",X"3F",X"57",X"08",X"CD",
		X"00",X"00",X"00",X"2D",X"D0",X"00",X"0D",X"2C",X"D0",X"0D",X"0D",X"D2",X"00",X"0C",X"53",X"FF",
		X"00",X"03",X"F2",X"FF",X"00",X"0D",X"D3",X"FF",X"00",X"0D",X"CF",X"FF",X"00",X"5F",X"DF",X"D7",
		X"00",X"FD",X"FF",X"2D",X"00",X"DD",X"FF",X"CD",X"D6",X"DF",X"FF",X"CD",X"DF",X"DF",X"5F",X"DF",
		X"DD",X"FF",X"76",X"FF",X"BD",X"FF",X"09",X"FF",X"2C",X"FF",X"09",X"DF",X"3F",X"57",X"08",X"BD",
		X"00",X"00",X"0D",X"32",X"00",X"00",X"03",X"D2",X"00",X"00",X"02",X"D3",X"00",X"00",X"53",X"FF",
		X"00",X"00",X"FD",X"DF",X"00",X"00",X"DD",X"3D",X"00",X"06",X"CD",X"FD",X"D0",X"5F",X"DF",X"5D",
		X"D0",X"FD",X"FF",X"DF",X"D0",X"DD",X"FF",X"FF",X"D6",X"DF",X"FF",X"FF",X"BF",X"DF",X"5F",X"FF",
		X"2D",X"FF",X"76",X"DF",X"3D",X"FF",X"09",X"BF",X"2D",X"FF",X"09",X"3C",X"CF",X"57",X"08",X"23",
		X"00",X"00",X"03",X"D3",X"00",X"00",X"00",X"DB",X"00",X"00",X"06",X"DD",X"00",X"00",X"5D",X"FF",
		X"00",X"00",X"FD",X"3F",X"00",X"00",X"DD",X"DF",X"00",X"06",X"CD",X"FF",X"D0",X"5D",X"DF",X"57",
		X"D0",X"FD",X"FF",X"FF",X"00",X"DD",X"FF",X"FF",X"26",X"DF",X"FF",X"FF",X"3F",X"DF",X"5F",X"FF",
		X"BD",X"FF",X"76",X"DF",X"DD",X"FF",X"09",X"2F",X"DD",X"FF",X"0D",X"33",X"DF",X"57",X"02",X"C2",
		X"FF",X"FF",X"00",X"DC",X"FF",X"FF",X"00",X"DC",X"FF",X"FF",X"06",X"2D",X"5F",X"FD",X"5F",X"FF",
		X"76",X"F3",X"FD",X"FF",X"09",X"F2",X"FD",X"FF",X"09",X"F3",X"D3",X"FF",X"D8",X"5D",X"DF",X"57",
		X"D0",X"FD",X"FF",X"44",X"00",X"DD",X"FF",X"44",X"06",X"DD",X"FF",X"44",X"5F",X"CF",X"54",X"44",
		X"FF",X"FF",X"76",X"44",X"FF",X"FF",X"09",X"44",X"DD",X"FF",X"09",X"44",X"CF",X"57",X"08",X"54",
		X"FF",X"FF",X"00",X"BD",X"FF",X"FF",X"00",X"2D",X"FF",X"F3",X"0D",X"2B",X"5F",X"F3",X"5D",X"FF",
		X"D6",X"F3",X"F3",X"FF",X"D9",X"F3",X"F3",X"FF",X"09",X"FB",X"CF",X"FF",X"08",X"5D",X"DF",X"57",
		X"00",X"FD",X"FF",X"44",X"00",X"D3",X"FF",X"44",X"06",X"D3",X"FF",X"44",X"5F",X"DF",X"54",X"44",
		X"DF",X"FF",X"76",X"44",X"DD",X"FF",X"09",X"44",X"CD",X"FF",X"09",X"44",X"3F",X"57",X"08",X"54",
		X"FF",X"FF",X"00",X"2D",X"DF",X"FF",X"0D",X"2C",X"DF",X"FD",X"0D",X"D2",X"5F",X"FC",X"53",X"FF",
		X"76",X"F3",X"F2",X"FF",X"09",X"FD",X"D3",X"FF",X"09",X"FD",X"CF",X"FF",X"08",X"5F",X"DF",X"57",
		X"00",X"FD",X"FF",X"44",X"00",X"DD",X"FF",X"44",X"D6",X"DF",X"FF",X"44",X"DF",X"DF",X"54",X"44",
		X"DD",X"FF",X"76",X"44",X"BD",X"FF",X"09",X"44",X"2C",X"FF",X"09",X"44",X"3F",X"57",X"08",X"54",
		X"FF",X"FF",X"0D",X"32",X"FF",X"FF",X"03",X"D2",X"FF",X"FF",X"02",X"D3",X"5F",X"FF",X"53",X"FF",
		X"76",X"FF",X"FD",X"FF",X"09",X"FF",X"DD",X"FF",X"09",X"FF",X"CD",X"FF",X"D8",X"5F",X"DF",X"57",
		X"D0",X"FD",X"FF",X"44",X"D0",X"DD",X"FF",X"44",X"D6",X"DF",X"FF",X"44",X"BF",X"DF",X"54",X"44",
		X"2D",X"FF",X"76",X"44",X"3D",X"FF",X"09",X"44",X"2D",X"FF",X"09",X"44",X"CF",X"57",X"08",X"54",
		X"FF",X"FF",X"03",X"D3",X"FF",X"FF",X"00",X"DB",X"FF",X"FF",X"06",X"DD",X"5F",X"FF",X"5D",X"FF",
		X"76",X"FF",X"FD",X"FF",X"09",X"FF",X"DD",X"FF",X"09",X"FF",X"CD",X"FF",X"D8",X"5D",X"DF",X"57",
		X"D0",X"FD",X"FF",X"44",X"00",X"DD",X"FF",X"44",X"26",X"DF",X"FF",X"44",X"3F",X"DF",X"54",X"44",
		X"BD",X"FF",X"76",X"44",X"DD",X"FF",X"09",X"44",X"DD",X"FF",X"09",X"44",X"DF",X"57",X"08",X"54",
		X"FF",X"FF",X"00",X"DC",X"FF",X"FF",X"00",X"DC",X"FF",X"FF",X"06",X"2D",X"5F",X"FD",X"5F",X"FF",
		X"76",X"F3",X"FD",X"FF",X"09",X"F2",X"FD",X"FF",X"09",X"F3",X"D3",X"FF",X"D8",X"5D",X"DF",X"57",
		X"D0",X"FD",X"FF",X"FF",X"00",X"DD",X"FF",X"FF",X"06",X"DD",X"FF",X"FF",X"5F",X"CF",X"5F",X"FF",
		X"FF",X"FF",X"76",X"FF",X"FF",X"FF",X"09",X"FF",X"DD",X"FF",X"09",X"FF",X"CF",X"57",X"08",X"5F",
		X"FF",X"FF",X"00",X"BD",X"FF",X"FF",X"00",X"2D",X"FF",X"F3",X"0D",X"2B",X"5F",X"F3",X"5D",X"FF",
		X"D6",X"F3",X"F3",X"FF",X"D9",X"F3",X"F3",X"FF",X"09",X"FB",X"CF",X"FF",X"08",X"5D",X"DF",X"57",
		X"00",X"FD",X"FF",X"FF",X"00",X"D3",X"FF",X"FF",X"06",X"D3",X"FF",X"FF",X"5F",X"DF",X"5F",X"FF",
		X"DF",X"FF",X"76",X"FF",X"DD",X"FF",X"09",X"FF",X"CD",X"FF",X"09",X"FF",X"3F",X"57",X"08",X"5F",
		X"FF",X"FF",X"00",X"2D",X"DF",X"FF",X"0D",X"2C",X"DF",X"FD",X"0D",X"D2",X"5F",X"FC",X"53",X"FF",
		X"76",X"F3",X"F2",X"FF",X"09",X"FD",X"D3",X"FF",X"09",X"FD",X"CF",X"FF",X"08",X"5F",X"DF",X"57",
		X"00",X"FD",X"FF",X"FF",X"00",X"DD",X"FF",X"FF",X"D6",X"DF",X"FF",X"FF",X"DF",X"DF",X"5F",X"FF",
		X"DD",X"FF",X"76",X"FF",X"BD",X"FF",X"09",X"FF",X"2C",X"FF",X"09",X"FF",X"3F",X"57",X"08",X"5F",
		X"FF",X"FF",X"0D",X"32",X"FF",X"FF",X"03",X"D2",X"FF",X"FF",X"02",X"D3",X"5F",X"FF",X"53",X"FF",
		X"76",X"FF",X"FD",X"FF",X"09",X"FF",X"DD",X"FF",X"09",X"FF",X"CD",X"FF",X"D8",X"5F",X"DF",X"57",
		X"D0",X"FD",X"FF",X"FF",X"D0",X"DD",X"FF",X"FF",X"D6",X"DF",X"FF",X"FF",X"BF",X"DF",X"5F",X"FF",
		X"2D",X"FF",X"76",X"FF",X"3D",X"FF",X"09",X"FF",X"2D",X"FF",X"09",X"FF",X"CF",X"57",X"08",X"5F",
		X"FF",X"FF",X"03",X"D3",X"FF",X"FF",X"00",X"DB",X"FF",X"FF",X"06",X"DD",X"5F",X"FF",X"5D",X"FF",
		X"76",X"FF",X"FD",X"FF",X"09",X"FF",X"DD",X"FF",X"09",X"FF",X"CD",X"FF",X"D8",X"5D",X"DF",X"57",
		X"D0",X"FD",X"FF",X"FF",X"00",X"DD",X"FF",X"FF",X"26",X"DF",X"FF",X"FF",X"3F",X"DF",X"5F",X"FF",
		X"BD",X"FF",X"76",X"FF",X"DD",X"FF",X"09",X"FF",X"DD",X"FF",X"09",X"FF",X"DF",X"57",X"08",X"5F",
		X"FF",X"FF",X"00",X"DC",X"FF",X"FF",X"00",X"DC",X"FF",X"FF",X"06",X"2D",X"5F",X"FD",X"5F",X"FF",
		X"76",X"F3",X"FD",X"DF",X"09",X"F2",X"FD",X"FF",X"09",X"F3",X"D3",X"FF",X"D8",X"5D",X"DF",X"57",
		X"D0",X"FD",X"FF",X"DF",X"00",X"DD",X"FF",X"DF",X"06",X"DD",X"FF",X"DF",X"5F",X"CF",X"5F",X"BF",
		X"FF",X"FF",X"76",X"3D",X"FF",X"FF",X"0D",X"2C",X"DD",X"FF",X"0D",X"33",X"CF",X"57",X"08",X"C3",
		X"FF",X"FF",X"00",X"BD",X"FF",X"FF",X"00",X"2D",X"FF",X"F3",X"0D",X"2B",X"5F",X"F3",X"5D",X"FF",
		X"D6",X"F3",X"F3",X"FF",X"D9",X"F3",X"F3",X"FF",X"09",X"FB",X"CF",X"FF",X"08",X"5D",X"DF",X"5D",
		X"00",X"FD",X"FF",X"DB",X"00",X"D3",X"FF",X"BD",X"06",X"D3",X"FF",X"2F",X"5F",X"DF",X"5D",X"2F",
		X"DF",X"FF",X"76",X"CF",X"DD",X"FF",X"09",X"DD",X"CD",X"FF",X"09",X"CD",X"3F",X"57",X"08",X"CD",
		X"FF",X"FF",X"00",X"2D",X"DF",X"FF",X"0D",X"2C",X"DF",X"FD",X"0D",X"D2",X"5F",X"FC",X"53",X"FF",
		X"76",X"F3",X"F2",X"FF",X"09",X"FD",X"D3",X"FF",X"09",X"FD",X"CF",X"FF",X"08",X"5F",X"DF",X"D7",
		X"00",X"FD",X"FF",X"2D",X"00",X"DD",X"FF",X"CD",X"D6",X"DF",X"FF",X"CD",X"DF",X"DF",X"5F",X"DF",
		X"DD",X"FF",X"76",X"FF",X"BD",X"FF",X"09",X"FF",X"2C",X"FF",X"09",X"DF",X"3F",X"57",X"08",X"BD",
		X"FF",X"FF",X"0D",X"32",X"FF",X"FF",X"03",X"D2",X"FF",X"FF",X"02",X"D3",X"5F",X"FF",X"53",X"FF",
		X"76",X"FF",X"FD",X"DF",X"09",X"FF",X"DD",X"3D",X"09",X"FF",X"CD",X"FD",X"D8",X"5F",X"DF",X"5D",
		X"D0",X"FD",X"FF",X"DF",X"D0",X"DD",X"FF",X"FF",X"D6",X"DF",X"FF",X"FF",X"BF",X"DF",X"5F",X"FF",
		X"2D",X"FF",X"76",X"DF",X"3D",X"FF",X"09",X"BF",X"2D",X"FF",X"09",X"3C",X"CF",X"57",X"08",X"23",
		X"FF",X"FF",X"03",X"D3",X"FF",X"FF",X"00",X"DB",X"FF",X"FF",X"06",X"DD",X"5F",X"FF",X"5D",X"FF",
		X"76",X"FF",X"FD",X"3F",X"09",X"FF",X"DD",X"DF",X"09",X"FF",X"CD",X"FF",X"D8",X"5D",X"DF",X"57",
		X"D0",X"FD",X"FF",X"FF",X"00",X"DD",X"FF",X"FF",X"26",X"DF",X"FF",X"FF",X"3F",X"DF",X"5F",X"FF",
		X"BD",X"FF",X"76",X"DF",X"DD",X"FF",X"09",X"2F",X"DD",X"FF",X"0D",X"33",X"DF",X"57",X"02",X"C2",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"06",X"FF",X"00",X"00",X"5F",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"06",X"FF",X"FF",X"00",X"5F",X"FF",X"57",
		X"00",X"FF",X"FF",X"44",X"00",X"FF",X"FF",X"44",X"06",X"FF",X"FF",X"44",X"5F",X"FF",X"54",X"44",
		X"FF",X"FF",X"76",X"44",X"FF",X"FF",X"09",X"44",X"FF",X"FF",X"09",X"44",X"FF",X"57",X"08",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"5F",
		X"00",X"00",X"00",X"6F",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"5F",
		X"00",X"00",X"00",X"6F",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"54",
		X"FF",X"44",X"00",X"44",X"FF",X"44",X"00",X"44",X"FF",X"44",X"06",X"44",X"54",X"44",X"54",X"44",
		X"76",X"44",X"44",X"44",X"09",X"44",X"44",X"44",X"09",X"44",X"44",X"44",X"08",X"54",X"44",X"57",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"06",X"44",X"44",X"44",X"54",X"44",X"54",X"44",
		X"44",X"44",X"76",X"44",X"44",X"44",X"09",X"44",X"44",X"44",X"09",X"44",X"44",X"57",X"08",X"54",
		X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"06",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"76",X"FF",X"FF",X"FF",X"09",X"FF",X"FF",X"FF",X"09",X"FF",X"FF",X"FF",X"08",X"5F",X"FF",X"57",
		X"00",X"FF",X"FF",X"44",X"00",X"FF",X"FF",X"44",X"06",X"FF",X"FF",X"44",X"5F",X"FF",X"54",X"44",
		X"FF",X"FF",X"76",X"44",X"FF",X"FF",X"09",X"44",X"FF",X"FF",X"09",X"44",X"FF",X"57",X"08",X"54",
		X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"06",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"76",X"FF",X"FF",X"FF",X"09",X"FF",X"FF",X"FF",X"09",X"FF",X"FF",X"FF",X"08",X"5F",X"FF",X"57",
		X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"06",X"FF",X"FF",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"FF",X"FF",X"76",X"FF",X"FF",X"FF",X"09",X"FF",X"FF",X"FF",X"09",X"FF",X"FF",X"57",X"08",X"5F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
