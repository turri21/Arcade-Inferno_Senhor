library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity inferno_bank_b is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of inferno_bank_b is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"20",X"49",X"4E",X"46",X"45",X"52",X"4E",X"4F",X"20",X"2D",X"20",X"43",X"4F",X"50",X"59",X"52",
		X"49",X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",X"38",X"34",X"20",X"57",X"49",
		X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",
		X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"00",X"02",X"00",X"00",X"02",X"00",X"00",X"A2",X"00",
		X"00",X"A2",X"00",X"00",X"22",X"00",X"0A",X"2D",X"00",X"0A",X"2D",X"00",X"A2",X"92",X"00",X"02",
		X"92",X"00",X"99",X"2D",X"00",X"02",X"2D",X"00",X"52",X"92",X"00",X"02",X"77",X"F0",X"79",X"2D",
		X"00",X"02",X"11",X"70",X"72",X"92",X"00",X"02",X"1A",X"70",X"1E",X"2D",X"00",X"02",X"F5",X"52",
		X"12",X"E2",X"00",X"0F",X"57",X"11",X"5E",X"ED",X"00",X"09",X"19",X"15",X"FE",X"20",X"00",X"05",
		X"10",X"17",X"02",X"00",X"00",X"00",X"FB",X"EA",X"F0",X"00",X"00",X"00",X"E1",X"5B",X"00",X"00",
		X"00",X"00",X"51",X"15",X"B0",X"00",X"00",X"00",X"BF",X"E1",X"50",X"00",X"00",X"00",X"70",X"71",
		X"50",X"00",X"00",X"00",X"7A",X"71",X"B0",X"00",X"00",X"00",X"7A",X"71",X"00",X"00",X"00",X"00",
		X"1A",X"77",X"00",X"00",X"00",X"00",X"1A",X"15",X"00",X"00",X"00",X"00",X"50",X"1A",X"00",X"00",
		X"00",X"00",X"70",X"59",X"00",X"00",X"00",X"00",X"10",X"15",X"00",X"00",X"00",X"00",X"10",X"15",
		X"00",X"00",X"00",X"00",X"50",X"1A",X"00",X"00",X"00",X"00",X"70",X"5B",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"07",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"50",
		X"00",X"01",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"D5",X"70",X"01",X"A7",X"00",X"00",X"55",
		X"99",X"9A",X"D0",X"02",X"51",X"F0",X"55",X"01",X"77",X"59",X"92",X"2D",X"00",X"03",X"25",X"17",
		X"11",X"15",X"E2",X"92",X"2D",X"00",X"00",X"00",X"29",X"19",X"15",X"FE",X"EE",X"2D",X"00",X"00",
		X"00",X"00",X"05",X"10",X"17",X"0E",X"EE",X"00",X"00",X"00",X"00",X"00",X"0D",X"FB",X"EA",X"FE",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"5B",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"51",X"15",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"E1",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"71",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7A",
		X"71",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7A",X"71",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1A",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"15",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"59",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"15",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",
		X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"5B",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"70",X"00",X"00",X"00",X"00",X"00",X"03",X"1A",X"70",
		X"00",X"00",X"00",X"00",X"00",X"E3",X"55",X"53",X"00",X"00",X"00",X"00",X"05",X"11",X"11",X"1E",
		X"E0",X"00",X"00",X"00",X"27",X"01",X"75",X"01",X"EE",X"00",X"00",X"0E",X"75",X"19",X"15",X"07",
		X"2E",X"E0",X"00",X"05",X"E5",X"10",X"17",X"FE",X"72",X"EF",X"00",X"05",X"2F",X"EE",X"AB",X"0D",
		X"5E",X"EF",X"00",X"09",X"E0",X"51",X"15",X"B0",X"35",X"EF",X"00",X"09",X"20",X"BF",X"E1",X"50",
		X"05",X"EF",X"00",X"09",X"E0",X"70",X"71",X"50",X"09",X"2F",X"00",X"09",X"E0",X"7A",X"71",X"B0",
		X"09",X"2F",X"00",X"0A",X"E0",X"7A",X"71",X"00",X"09",X"20",X"00",X"00",X"D0",X"1A",X"77",X"00",
		X"09",X"D0",X"00",X"00",X"00",X"1A",X"15",X"00",X"0A",X"00",X"00",X"00",X"00",X"50",X"1A",X"00",
		X"0D",X"00",X"00",X"00",X"00",X"70",X"59",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"15",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"1A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"5B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"20",X"00",X"00",X"0A",X"20",X"00",X"0A",X"20",X"00",
		X"00",X"02",X"20",X"00",X"A2",X"D0",X"00",X"00",X"A2",X"D0",X"0A",X"29",X"20",X"00",X"00",X"29",
		X"20",X"09",X"92",X"D0",X"00",X"00",X"22",X"D0",X"05",X"29",X"20",X"00",X"00",X"27",X"7F",X"07",
		X"92",X"D0",X"00",X"00",X"21",X"17",X"07",X"29",X"20",X"00",X"00",X"21",X"A7",X"01",X"E2",X"D0",
		X"00",X"00",X"2F",X"55",X"21",X"2E",X"20",X"00",X"00",X"F5",X"71",X"15",X"EE",X"D0",X"00",X"00",
		X"91",X"91",X"5F",X"E2",X"00",X"00",X"00",X"51",X"01",X"70",X"20",X"00",X"00",X"00",X"0F",X"BE",
		X"AF",X"00",X"00",X"00",X"00",X"0E",X"15",X"B0",X"00",X"00",X"00",X"00",X"05",X"11",X"5B",X"00",
		X"00",X"00",X"00",X"0B",X"FE",X"15",X"00",X"00",X"00",X"00",X"07",X"70",X"15",X"A0",X"00",X"00",
		X"00",X"05",X"70",X"1B",X"50",X"00",X"00",X"00",X"09",X"70",X"71",X"90",X"00",X"00",X"00",X"00",
		X"19",X"51",X"70",X"00",X"00",X"00",X"00",X"01",X"07",X"1A",X"00",X"00",X"00",X"00",X"00",X"70",
		X"55",X"50",X"00",X"00",X"00",X"00",X"01",X"01",X"5A",X"00",X"00",X"00",X"00",X"00",X"70",X"15",
		X"00",X"00",X"00",X"00",X"00",X"05",X"01",X"90",X"00",X"00",X"00",X"00",X"00",X"90",X"79",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"77",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"11",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"57",X"00",X"1A",X"70",X"00",X"05",X"59",X"99",X"AD",X"00",X"00",X"00",X"25",X"1F",X"05",X"50",
		X"17",X"75",X"99",X"22",X"D0",X"00",X"00",X"00",X"32",X"51",X"71",X"11",X"5E",X"29",X"22",X"D0",
		X"00",X"00",X"00",X"00",X"02",X"91",X"91",X"5F",X"EE",X"E2",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"51",X"01",X"70",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"BE",X"0F",
		X"ED",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"B1",X"70",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"51",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"51",X"11",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"51",X"77",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"11",
		X"51",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"51",X"70",X"00",
		X"00",X"07",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"17",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"A7",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"35",X"55",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"59",X"71",X"11",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"91",X"91",X"50",X"1E",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"51",X"01",X"70",X"72",X"EE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"9E",X"2E",X"CA",X"EE",X"E7",X"2E",X"F9",X"00",X"00",X"00",X"00",X"00",X"92",
		X"EE",X"0A",X"E5",X"D5",X"EE",X"F1",X"77",X"50",X"00",X"00",X"00",X"9E",X"E0",X"00",X"04",X"53",
		X"5E",X"F1",X"15",X"11",X"51",X"90",X"00",X"92",X"E0",X"00",X"00",X"00",X"5E",X"F0",X"00",X"00",
		X"09",X"51",X"70",X"9E",X"E0",X"00",X"00",X"00",X"92",X"F0",X"00",X"00",X"00",X"00",X"00",X"AE",
		X"F0",X"00",X"00",X"00",X"92",X"F0",X"00",X"00",X"00",X"00",X"00",X"AE",X"00",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"02",X"00",
		X"00",X"02",X"A0",X"00",X"02",X"A0",X"00",X"0D",X"2A",X"00",X"02",X"20",X"00",X"02",X"92",X"A0",
		X"0D",X"2A",X"00",X"0D",X"29",X"90",X"02",X"92",X"00",X"02",X"92",X"50",X"0D",X"22",X"00",X"0D",
		X"29",X"70",X"F7",X"72",X"00",X"02",X"92",X"70",X"71",X"12",X"00",X"0D",X"2E",X"10",X"7A",X"12",
		X"00",X"02",X"E2",X"12",X"55",X"F2",X"00",X"0D",X"EE",X"51",X"17",X"5F",X"00",X"00",X"2E",X"F5",
		X"19",X"19",X"00",X"00",X"02",X"07",X"10",X"15",X"00",X"00",X"00",X"FA",X"EB",X"F0",X"00",X"00",
		X"00",X"0B",X"51",X"E0",X"00",X"00",X"00",X"B5",X"11",X"50",X"00",X"00",X"00",X"51",X"EF",X"B0",
		X"00",X"00",X"00",X"51",X"70",X"70",X"00",X"00",X"00",X"B1",X"7A",X"70",X"00",X"00",X"00",X"01",
		X"7A",X"70",X"00",X"00",X"00",X"07",X"7A",X"10",X"00",X"00",X"00",X"05",X"1A",X"10",X"00",X"00",
		X"00",X"0A",X"10",X"50",X"00",X"00",X"00",X"09",X"50",X"70",X"00",X"00",X"00",X"05",X"10",X"10",
		X"00",X"00",X"00",X"05",X"10",X"10",X"00",X"00",X"00",X"0A",X"10",X"50",X"00",X"00",X"00",X"0B",
		X"50",X"70",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"11",X"00",X"00",X"50",X"DA",X"99",X"95",
		X"50",X"00",X"07",X"A1",X"00",X"75",X"D0",X"0D",X"22",X"99",X"57",X"71",X"05",X"50",X"F1",X"52",
		X"00",X"00",X"0D",X"22",X"92",X"E5",X"11",X"17",X"15",X"23",X"00",X"00",X"00",X"0D",X"2E",X"EE",
		X"F5",X"19",X"19",X"20",X"00",X"00",X"00",X"00",X"0E",X"EE",X"07",X"10",X"15",X"00",X"00",X"00",
		X"00",X"00",X"00",X"DE",X"FA",X"EB",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0B",X"51",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B5",X"11",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"51",X"EF",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"51",X"70",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B1",X"7A",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"7A",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"7A",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"1A",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"10",
		X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"50",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"10",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"50",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F7",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"7A",X"13",X"00",X"00",X"00",X"00",X"00",X"03",X"55",X"53",X"E0",X"00",X"00",X"00",
		X"00",X"EE",X"11",X"11",X"15",X"00",X"00",X"00",X"0E",X"E1",X"05",X"71",X"07",X"20",X"00",X"00",
		X"EE",X"27",X"05",X"19",X"15",X"7E",X"00",X"0F",X"E2",X"7E",X"F7",X"10",X"15",X"E5",X"00",X"0F",
		X"EE",X"5D",X"0B",X"AE",X"EF",X"25",X"00",X"0F",X"E5",X"30",X"B5",X"11",X"50",X"E9",X"00",X"0F",
		X"E5",X"00",X"51",X"EF",X"B0",X"29",X"00",X"0F",X"29",X"00",X"51",X"70",X"70",X"E9",X"00",X"0F",
		X"29",X"00",X"B1",X"7A",X"70",X"E9",X"00",X"00",X"29",X"00",X"01",X"7A",X"70",X"EA",X"00",X"00",
		X"D9",X"00",X"07",X"7A",X"10",X"D0",X"00",X"00",X"0A",X"00",X"05",X"1A",X"10",X"00",X"00",X"00",
		X"0D",X"00",X"0A",X"10",X"50",X"00",X"00",X"00",X"00",X"00",X"09",X"50",X"70",X"00",X"00",X"00",
		X"00",X"00",X"05",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"05",X"10",X"10",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"10",X"50",X"00",X"00",X"00",X"00",X"00",X"0B",X"50",X"70",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"20",X"00",X"00",X"00",
		X"2A",X"00",X"00",X"2A",X"00",X"00",X"00",X"D2",X"A0",X"00",X"22",X"00",X"00",X"00",X"29",X"2A",
		X"00",X"D2",X"A0",X"00",X"00",X"D2",X"99",X"00",X"29",X"20",X"00",X"00",X"29",X"25",X"00",X"D2",
		X"20",X"00",X"00",X"D2",X"97",X"0F",X"77",X"20",X"00",X"00",X"29",X"27",X"07",X"11",X"20",X"00",
		X"00",X"D2",X"E1",X"07",X"A1",X"20",X"00",X"00",X"2E",X"21",X"25",X"5F",X"20",X"00",X"00",X"DE",
		X"E5",X"11",X"75",X"F0",X"00",X"00",X"02",X"EF",X"51",X"91",X"90",X"00",X"00",X"00",X"20",X"71",
		X"01",X"50",X"00",X"00",X"00",X"0F",X"AE",X"BF",X"00",X"00",X"00",X"00",X"00",X"B5",X"1E",X"00",
		X"00",X"00",X"00",X"0B",X"51",X"15",X"00",X"00",X"00",X"00",X"05",X"1E",X"FB",X"00",X"00",X"00",
		X"00",X"A5",X"10",X"77",X"00",X"00",X"00",X"00",X"5B",X"10",X"75",X"00",X"00",X"00",X"00",X"91",
		X"70",X"79",X"00",X"00",X"00",X"00",X"71",X"59",X"10",X"00",X"00",X"00",X"0A",X"17",X"01",X"00",
		X"00",X"00",X"00",X"55",X"50",X"70",X"00",X"00",X"00",X"0A",X"51",X"01",X"00",X"00",X"00",X"00",
		X"05",X"10",X"70",X"00",X"00",X"00",X"00",X"91",X"05",X"00",X"00",X"00",X"00",X"09",X"70",X"90",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F7",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"10",
		X"00",X"05",X"00",X"00",X"0D",X"A9",X"99",X"55",X"00",X"00",X"7A",X"10",X"07",X"5D",X"00",X"00",
		X"00",X"D2",X"29",X"95",X"77",X"10",X"55",X"0F",X"15",X"20",X"00",X"00",X"00",X"00",X"D2",X"29",
		X"2E",X"51",X"11",X"71",X"52",X"30",X"00",X"00",X"00",X"00",X"00",X"D2",X"EE",X"EF",X"51",X"91",
		X"92",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"E0",X"71",X"01",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0D",X"EF",X"0E",X"B0",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"71",X"B5",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"11",X"51",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"11",X"11",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"57",X"71",X"59",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"91",X"51",X"15",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"77",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"A1",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"35",X"55",
		X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"E1",X"11",X"79",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"10",X"51",X"91",X"95",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"E2",X"70",X"71",X"01",X"59",X"90",X"00",X"00",X"00",X"00",X"09",X"FE",X"27",X"EE",X"EA",
		X"CE",X"2E",X"90",X"00",X"00",X"00",X"57",X"71",X"FE",X"E5",X"D5",X"EA",X"0E",X"E2",X"90",X"00",
		X"91",X"51",X"15",X"11",X"FE",X"53",X"54",X"00",X"00",X"EE",X"90",X"71",X"59",X"00",X"00",X"00",
		X"FE",X"50",X"00",X"00",X"00",X"E2",X"90",X"00",X"00",X"00",X"00",X"00",X"F2",X"90",X"00",X"00",
		X"00",X"EE",X"90",X"00",X"00",X"00",X"00",X"00",X"F2",X"90",X"00",X"00",X"00",X"FE",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"02",X"90",X"00",X"00",X"00",X"0E",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"90",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0D",X"E9",X"99",X"55",X"50",X"00",X"00",X"01",X"A7",X"00",X"00",X"55",X"99",X"9A",X"D0",
		X"00",X"00",X"00",X"DD",X"22",X"99",X"55",X"77",X"10",X"00",X"55",X"01",X"77",X"59",X"92",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"0D",X"22",X"92",X"E9",X"21",X"17",X"79",X"15",X"E2",X"92",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"2E",X"E2",X"E2",X"11",X"17",X"5E",X"EE",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"EE",X"2E",X"E9",X"77",X"0E",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DE",X"E7",X"11",X"1E",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"11",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"1E",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"11",X"11",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"95",X"17",X"75",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"51",X"15",X"19",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"17",X"00",X"00",X"00",X"07",
		X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"17",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"A7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"35",X"55",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D1",X"71",
		X"19",X"1E",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"11",X"11",X"19",X"9E",X"E5",X"00",
		X"00",X"00",X"00",X"00",X"00",X"95",X"5E",X"E9",X"75",X"17",X"15",X"00",X"00",X"00",X"00",X"00",
		X"00",X"59",X"2E",X"EE",X"11",X"11",X"11",X"59",X"00",X"00",X"00",X"00",X"00",X"52",X"EE",X"ED",
		X"05",X"11",X"11",X"11",X"77",X"50",X"00",X"00",X"00",X"5E",X"E2",X"D0",X"00",X"05",X"11",X"11",
		X"15",X"11",X"51",X"90",X"00",X"92",X"EE",X"00",X"00",X"00",X"5E",X"F0",X"00",X"00",X"09",X"51",
		X"70",X"92",X"2D",X"00",X"00",X"00",X"92",X"D0",X"00",X"00",X"00",X"00",X"00",X"A2",X"20",X"00",
		X"00",X"00",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"AE",X"E0",X"00",X"00",X"00",X"9D",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"D0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DA",X"99",X"95",
		X"50",X"00",X"07",X"A1",X"00",X"00",X"00",X"55",X"59",X"99",X"ED",X"00",X"00",X"00",X"0D",X"22",
		X"99",X"57",X"71",X"05",X"50",X"00",X"17",X"75",X"59",X"92",X"2D",X"D0",X"00",X"00",X"00",X"00",
		X"0D",X"22",X"92",X"E5",X"19",X"77",X"11",X"29",X"E2",X"92",X"2D",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"2E",X"EE",X"57",X"11",X"12",X"E2",X"EE",X"2D",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"EE",X"07",X"79",X"EE",X"2E",X"ED",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"DE",X"11",X"17",X"EE",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"11",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"11",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"11",X"15",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"77",X"15",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"15",X"11",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"A1",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"35",X"55",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5E",X"19",X"11",
		X"71",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"EE",X"99",X"11",X"11",X"15",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"17",X"15",X"79",X"EE",X"55",X"90",X"00",X"00",X"00",X"00",X"09",
		X"51",X"11",X"11",X"1E",X"EE",X"29",X"50",X"00",X"00",X"00",X"57",X"71",X"11",X"11",X"15",X"0D",
		X"EE",X"E2",X"50",X"00",X"91",X"51",X"15",X"11",X"11",X"15",X"00",X"00",X"D2",X"EE",X"50",X"71",
		X"59",X"00",X"00",X"00",X"FE",X"50",X"00",X"00",X"0E",X"E2",X"90",X"00",X"00",X"00",X"00",X"00",
		X"D2",X"90",X"00",X"00",X"0D",X"22",X"90",X"00",X"00",X"00",X"00",X"00",X"0A",X"90",X"00",X"00",
		X"00",X"22",X"A0",X"00",X"00",X"00",X"00",X"00",X"0D",X"90",X"00",X"00",X"00",X"EE",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"D2",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"09",X"55",X"55",X"59",X"00",
		X"00",X"00",X"05",X"5A",X"55",X"55",X"00",X"00",X"00",X"05",X"50",X"05",X"5A",X"00",X"00",X"00",
		X"05",X"50",X"05",X"50",X"00",X"00",X"00",X"09",X"50",X"05",X"50",X"00",X"00",X"00",X"00",X"55",
		X"09",X"5A",X"00",X"00",X"00",X"00",X"55",X"00",X"55",X"00",X"00",X"00",X"05",X"55",X"00",X"55",
		X"00",X"00",X"08",X"55",X"A8",X"88",X"55",X"88",X"00",X"00",X"88",X"88",X"A5",X"55",X"88",X"80",
		X"00",X"88",X"88",X"55",X"A8",X"88",X"00",X"00",X"00",X"88",X"88",X"88",X"80",X"00",X"00",X"55",
		X"55",X"50",X"00",X"00",X"09",X"85",X"55",X"50",X"00",X"00",X"0A",X"55",X"59",X"00",X"00",X"00",
		X"09",X"55",X"00",X"00",X"00",X"00",X"05",X"50",X"00",X"00",X"00",X"00",X"05",X"59",X"00",X"00",
		X"00",X"00",X"0A",X"95",X"50",X"00",X"00",X"00",X"00",X"A9",X"59",X"88",X"80",X"00",X"05",X"98",
		X"55",X"88",X"88",X"00",X"55",X"A9",X"5A",X"88",X"80",X"00",X"00",X"05",X"58",X"88",X"00",X"00",
		X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"55",X"55",X"50",
		X"00",X"00",X"00",X"98",X"55",X"90",X"00",X"00",X"00",X"A9",X"55",X"00",X"00",X"00",X"00",X"A5",
		X"59",X"00",X"00",X"00",X"00",X"05",X"5A",X"5A",X"00",X"00",X"00",X"05",X"9A",X"95",X"5A",X"00",
		X"00",X"09",X"50",X"8A",X"59",X"00",X"00",X"05",X"90",X"0A",X"58",X"00",X"00",X"05",X"50",X"8A",
		X"58",X"80",X"00",X"05",X"58",X"88",X"88",X"80",X"00",X"95",X"58",X"88",X"88",X"00",X"05",X"55",
		X"88",X"80",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"05",X"55",X"55",X"59",
		X"00",X"00",X"00",X"55",X"5A",X"55",X"55",X"00",X"00",X"05",X"59",X"00",X"05",X"5A",X"00",X"00",
		X"95",X"50",X"00",X"05",X"50",X"00",X"00",X"A5",X"55",X"90",X"09",X"50",X"00",X"00",X"00",X"A5",
		X"50",X"0A",X"55",X"00",X"00",X"00",X"05",X"90",X"00",X"55",X"00",X"00",X"00",X"05",X"00",X"00",
		X"55",X"00",X"00",X"08",X"88",X"88",X"A5",X"55",X"80",X"00",X"00",X"08",X"88",X"55",X"A8",X"88",
		X"00",X"00",X"00",X"08",X"88",X"88",X"80",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",
		X"00",X"00",X"05",X"55",X"55",X"59",X"00",X"00",X"00",X"00",X"55",X"5A",X"55",X"59",X"00",X"00",
		X"00",X"0A",X"55",X"00",X"95",X"5A",X"00",X"00",X"00",X"05",X"50",X"00",X"05",X"50",X"00",X"00",
		X"00",X"05",X"A0",X"00",X"05",X"5A",X"9A",X"00",X"00",X"05",X"90",X"00",X"09",X"59",X"95",X"00",
		X"00",X"05",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"05",X"50",X"00",X"00",X"00",X"5A",X"00",
		X"0A",X"55",X"58",X"88",X"88",X"88",X"88",X"00",X"05",X"5A",X"88",X"88",X"88",X"88",X"00",X"00",
		X"00",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"09",
		X"8A",X"55",X"50",X"00",X"00",X"00",X"A9",X"A5",X"59",X"00",X"00",X"00",X"00",X"9A",X"95",X"58",
		X"00",X"00",X"00",X"00",X"AA",X"55",X"AA",X"A0",X"00",X"00",X"00",X"00",X"55",X"A9",X"58",X"00",
		X"00",X"00",X"00",X"55",X"89",X"88",X"80",X"00",X"00",X"00",X"A5",X"50",X"88",X"88",X"80",X"00",
		X"00",X"00",X"55",X"00",X"88",X"88",X"00",X"00",X"00",X"05",X"58",X"88",X"80",X"00",X"00",X"00",
		X"A5",X"98",X"88",X"80",X"00",X"00",X"00",X"55",X"88",X"88",X"80",X"00",X"00",X"55",X"55",X"50",
		X"00",X"09",X"85",X"55",X"50",X"00",X"09",X"55",X"5A",X"00",X"00",X"95",X"59",X"00",X"00",X"00",
		X"55",X"AA",X"95",X"A0",X"00",X"99",X"55",X"55",X"90",X"00",X"09",X"A0",X"09",X"50",X"00",X"05",
		X"58",X"8A",X"90",X"00",X"05",X"58",X"88",X"00",X"00",X"A5",X"58",X"88",X"88",X"00",X"55",X"A8",
		X"88",X"88",X"80",X"08",X"88",X"88",X"88",X"00",X"00",X"00",X"09",X"11",X"15",X"D0",X"00",X"00",
		X"00",X"97",X"77",X"77",X"90",X"00",X"00",X"00",X"98",X"88",X"87",X"90",X"00",X"00",X"00",X"A8",
		X"98",X"89",X"A0",X"00",X"00",X"00",X"A8",X"A8",X"88",X"5D",X"00",X"00",X"05",X"A8",X"88",X"A5",
		X"55",X"00",X"00",X"5A",X"8A",X"A9",X"55",X"59",X"00",X"05",X"A8",X"8A",X"55",X"5A",X"AA",X"00",
		X"A7",X"85",X"95",X"5A",X"A9",X"90",X"00",X"1E",X"55",X"5A",X"A9",X"59",X"00",X"00",X"00",X"00",
		X"95",X"55",X"50",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"50",X"00",X"00",X"00",X"00",X"09",X"18",X"50",X"00",X"00",
		X"00",X"00",X"05",X"87",X"55",X"00",X"00",X"00",X"00",X"95",X"58",X"95",X"50",X"00",X"00",X"05",
		X"58",X"88",X"88",X"55",X"00",X"00",X"95",X"89",X"11",X"15",X"D5",X"90",X"00",X"58",X"97",X"77",
		X"77",X"99",X"5A",X"00",X"58",X"58",X"88",X"87",X"98",X"5A",X"00",X"9A",X"A8",X"98",X"85",X"A8",
		X"5A",X"00",X"A5",X"A8",X"A8",X"8A",X"A5",X"5A",X"00",X"09",X"A8",X"88",X"88",X"55",X"90",X"00",
		X"0A",X"5A",X"8A",X"A5",X"99",X"00",X"00",X"00",X"55",X"A5",X"55",X"AA",X"00",X"00",X"00",X"55",
		X"95",X"59",X"A0",X"00",X"00",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"95",X"55",X"50",
		X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"09",X"55",X"55",X"59",X"00",
		X"00",X"00",X"05",X"55",X"5A",X"55",X"00",X"00",X"00",X"0A",X"55",X"00",X"55",X"00",X"00",X"00",
		X"00",X"55",X"00",X"55",X"00",X"00",X"00",X"00",X"55",X"00",X"59",X"00",X"00",X"00",X"0A",X"59",
		X"05",X"50",X"00",X"00",X"00",X"05",X"50",X"05",X"50",X"00",X"00",X"00",X"05",X"50",X"05",X"55",
		X"00",X"00",X"08",X"85",X"58",X"88",X"A5",X"58",X"00",X"88",X"85",X"55",X"A8",X"88",X"80",X"00",
		X"08",X"88",X"A5",X"58",X"88",X"80",X"00",X"00",X"88",X"88",X"88",X"80",X"00",X"00",X"00",X"00",
		X"55",X"55",X"50",X"00",X"00",X"00",X"55",X"55",X"89",X"00",X"00",X"00",X"09",X"55",X"5A",X"00",
		X"00",X"00",X"00",X"05",X"59",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"09",
		X"55",X"00",X"00",X"00",X"00",X"55",X"9A",X"00",X"00",X"88",X"89",X"59",X"A0",X"00",X"08",X"88",
		X"85",X"58",X"95",X"00",X"00",X"88",X"8A",X"59",X"A5",X"50",X"00",X"08",X"88",X"55",X"00",X"00",
		X"00",X"00",X"08",X"80",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"55",X"55",
		X"50",X"00",X"00",X"00",X"95",X"58",X"90",X"00",X"00",X"00",X"05",X"59",X"A0",X"00",X"00",X"00",
		X"09",X"55",X"A0",X"00",X"00",X"0A",X"5A",X"55",X"00",X"00",X"0A",X"55",X"9A",X"95",X"00",X"00",
		X"09",X"5A",X"80",X"59",X"00",X"00",X"08",X"5A",X"00",X"95",X"00",X"00",X"88",X"5A",X"80",X"55",
		X"00",X"00",X"88",X"88",X"88",X"55",X"00",X"00",X"08",X"88",X"88",X"55",X"90",X"00",X"00",X"00",
		X"88",X"85",X"55",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"09",X"55",X"55",X"55",
		X"00",X"00",X"00",X"05",X"55",X"5A",X"55",X"50",X"00",X"00",X"0A",X"55",X"00",X"09",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"55",X"90",X"00",X"00",X"59",X"00",X"95",X"55",X"A0",X"00",X"05",
		X"5A",X"00",X"55",X"A0",X"00",X"00",X"05",X"50",X"00",X"95",X"00",X"00",X"00",X"05",X"50",X"00",
		X"05",X"00",X"00",X"00",X"85",X"55",X"A8",X"88",X"88",X"00",X"08",X"88",X"A5",X"58",X"88",X"00",
		X"00",X"00",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"00",
		X"00",X"09",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"09",X"55",X"5A",X"55",X"50",X"00",X"00",
		X"00",X"0A",X"55",X"90",X"05",X"5A",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"55",X"00",X"00",
		X"0A",X"9A",X"55",X"00",X"00",X"A5",X"00",X"00",X"05",X"99",X"59",X"00",X"00",X"95",X"00",X"00",
		X"05",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"0A",X"50",X"00",X"00",X"00",X"55",X"00",X"00",
		X"08",X"88",X"88",X"88",X"88",X"55",X"5A",X"00",X"00",X"08",X"88",X"88",X"88",X"8A",X"55",X"00",
		X"00",X"00",X"00",X"08",X"88",X"88",X"80",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",
		X"00",X"00",X"55",X"5A",X"89",X"00",X"00",X"00",X"00",X"09",X"55",X"A9",X"A0",X"00",X"00",X"00",
		X"08",X"55",X"9A",X"90",X"00",X"00",X"00",X"AA",X"A5",X"5A",X"A0",X"00",X"00",X"08",X"59",X"A5",
		X"50",X"00",X"00",X"00",X"88",X"89",X"85",X"50",X"00",X"00",X"88",X"88",X"80",X"55",X"A0",X"00",
		X"08",X"88",X"80",X"05",X"50",X"00",X"00",X"00",X"88",X"88",X"55",X"00",X"00",X"00",X"00",X"88",
		X"88",X"95",X"A0",X"00",X"00",X"00",X"88",X"88",X"85",X"50",X"00",X"00",X"00",X"55",X"55",X"50",
		X"00",X"00",X"55",X"55",X"89",X"00",X"00",X"0A",X"55",X"59",X"00",X"00",X"00",X"09",X"55",X"90",
		X"00",X"A5",X"9A",X"A5",X"50",X"00",X"95",X"55",X"59",X"90",X"00",X"59",X"00",X"A9",X"00",X"00",
		X"9A",X"88",X"55",X"00",X"00",X"08",X"88",X"55",X"00",X"08",X"88",X"88",X"55",X"A0",X"88",X"88",
		X"88",X"A5",X"50",X"08",X"88",X"88",X"88",X"00",X"00",X"D5",X"11",X"19",X"00",X"00",X"00",X"00",
		X"97",X"77",X"77",X"90",X"00",X"00",X"00",X"97",X"88",X"88",X"90",X"00",X"00",X"00",X"A9",X"88",
		X"98",X"A0",X"00",X"00",X"0D",X"58",X"88",X"A8",X"A0",X"00",X"00",X"05",X"55",X"A8",X"88",X"A5",
		X"00",X"00",X"09",X"55",X"59",X"AA",X"8A",X"50",X"00",X"0A",X"AA",X"55",X"5A",X"88",X"A5",X"00",
		X"00",X"99",X"AA",X"55",X"95",X"87",X"A0",X"00",X"09",X"59",X"AA",X"55",X"5E",X"10",X"00",X"00",
		X"55",X"55",X"90",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"00",X"00",X"00",X"00",X"00",X"00",X"58",X"19",X"00",
		X"00",X"00",X"00",X"05",X"57",X"85",X"00",X"00",X"00",X"00",X"55",X"98",X"55",X"90",X"00",X"00",
		X"05",X"58",X"88",X"88",X"55",X"00",X"00",X"95",X"D5",X"11",X"19",X"85",X"90",X"0A",X"59",X"97",
		X"77",X"77",X"98",X"50",X"0A",X"58",X"97",X"88",X"88",X"58",X"50",X"0A",X"58",X"A5",X"88",X"98",
		X"AA",X"90",X"0A",X"55",X"AA",X"88",X"A8",X"A5",X"A0",X"00",X"95",X"58",X"88",X"88",X"A9",X"00",
		X"00",X"09",X"95",X"AA",X"8A",X"5A",X"00",X"00",X"0A",X"A5",X"55",X"A5",X"50",X"00",X"00",X"00",
		X"A9",X"55",X"95",X"50",X"00",X"00",X"00",X"09",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"55",
		X"55",X"90",X"00",X"00",X"55",X"55",X"50",X"00",X"09",X"55",X"59",X"90",X"00",X"05",X"55",X"AA",
		X"90",X"00",X"05",X"50",X"A9",X"A0",X"00",X"05",X"50",X"05",X"A0",X"00",X"05",X"50",X"09",X"50",
		X"00",X"09",X"50",X"0A",X"5A",X"00",X"00",X"5A",X"80",X"59",X"00",X"00",X"59",X"85",X"55",X"00",
		X"5A",X"55",X"88",X"59",X"80",X"95",X"59",X"88",X"88",X"80",X"00",X"5A",X"88",X"88",X"00",X"00",
		X"08",X"88",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"95",X"55",X"59",X"90",X"00",
		X"05",X"55",X"5A",X"AA",X"90",X"00",X"A5",X"50",X"00",X"A9",X"A0",X"00",X"09",X"59",X"00",X"05",
		X"A0",X"00",X"00",X"59",X"00",X"05",X"90",X"00",X"00",X"95",X"A0",X"09",X"50",X"00",X"00",X"54",
		X"A0",X"00",X"5A",X"00",X"05",X"4A",X"00",X"00",X"59",X"00",X"09",X"A0",X"00",X"95",X"55",X"00",
		X"00",X"00",X"08",X"88",X"5A",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"08",X"88",X"88",
		X"80",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"59",
		X"90",X"00",X"00",X"00",X"00",X"00",X"55",X"59",X"AA",X"90",X"00",X"00",X"00",X"00",X"09",X"59",
		X"A0",X"A9",X"A0",X"00",X"00",X"00",X"00",X"05",X"9A",X"00",X"A5",X"90",X"00",X"00",X"00",X"00",
		X"05",X"50",X"00",X"05",X"5A",X"00",X"00",X"00",X"0A",X"05",X"50",X"00",X"0A",X"55",X"99",X"D0",
		X"00",X"05",X"95",X"90",X"00",X"00",X"00",X"54",X"A0",X"00",X"00",X"55",X"A0",X"00",X"00",X"00",
		X"54",X"00",X"00",X"00",X"05",X"08",X"88",X"88",X"85",X"94",X"88",X"00",X"00",X"00",X"08",X"88",
		X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"80",X"00",X"00",X"00",X"55",
		X"55",X"50",X"00",X"09",X"55",X"59",X"90",X"00",X"05",X"55",X"AA",X"90",X"00",X"05",X"5A",X"8A",
		X"A0",X"00",X"05",X"58",X"AA",X"9A",X"00",X"09",X"58",X"A9",X"4A",X"00",X"0A",X"59",X"05",X"4A",
		X"00",X"00",X"55",X"09",X"50",X"00",X"00",X"55",X"88",X"80",X"00",X"55",X"55",X"88",X"88",X"00",
		X"05",X"59",X"88",X"88",X"00",X"00",X"5A",X"88",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",
		X"A5",X"55",X"59",X"90",X"0A",X"55",X"55",X"AA",X"90",X"A5",X"59",X"AA",X"A9",X"A0",X"95",X"9A",
		X"8A",X"9A",X"00",X"A5",X"55",X"55",X"90",X"00",X"00",X"09",X"54",X"50",X"00",X"00",X"00",X"54",
		X"50",X"00",X"00",X"00",X"59",X"AA",X"00",X"00",X"00",X"0A",X"A9",X"00",X"00",X"00",X"A5",X"9A",
		X"00",X"00",X"88",X"55",X"A8",X"00",X"08",X"88",X"88",X"88",X"80",X"08",X"88",X"88",X"80",X"00",
		X"00",X"88",X"80",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"55",X"55",X"59",
		X"00",X"00",X"95",X"55",X"59",X"99",X"00",X"A5",X"55",X"59",X"AA",X"9A",X"00",X"95",X"5A",X"00",
		X"AA",X"A0",X"00",X"95",X"A0",X"0A",X"9A",X"00",X"00",X"05",X"90",X"09",X"A0",X"00",X"00",X"09",
		X"50",X"09",X"59",X"00",X"00",X"55",X"50",X"00",X"95",X"50",X"00",X"A9",X"50",X"00",X"0A",X"5A",
		X"00",X"00",X"00",X"88",X"89",X"30",X"00",X"00",X"88",X"88",X"85",X"A0",X"00",X"88",X"88",X"88",
		X"88",X"80",X"00",X"00",X"08",X"88",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"0A",X"55",
		X"55",X"50",X"00",X"AA",X"55",X"59",X"90",X"00",X"AA",X"55",X"9A",X"00",X"00",X"0A",X"55",X"A0",
		X"00",X"00",X"00",X"95",X"88",X"00",X"00",X"08",X"A5",X"5A",X"00",X"00",X"08",X"88",X"55",X"A0",
		X"00",X"00",X"88",X"85",X"5A",X"00",X"00",X"00",X"89",X"55",X"00",X"00",X"00",X"55",X"9A",X"00",
		X"00",X"08",X"88",X"80",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"07",X"11",X"1E",X"00",
		X"00",X"1E",X"F0",X"71",X"17",X"75",X"00",X"00",X"89",X"78",X"89",X"77",X"59",X"00",X"00",X"05",
		X"98",X"88",X"55",X"59",X"A0",X"00",X"0A",X"58",X"88",X"99",X"9F",X"A9",X"00",X"09",X"55",X"8F",
		X"FF",X"FA",X"95",X"00",X"0A",X"55",X"55",X"55",X"99",X"59",X"00",X"00",X"A9",X"55",X"55",X"99",
		X"9A",X"00",X"00",X"00",X"A9",X"99",X"9A",X"90",X"00",X"00",X"00",X"A5",X"99",X"A5",X"00",X"00",
		X"00",X"00",X"55",X"5A",X"50",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"09",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"95",X"78",X"50",X"00",X"00",X"00",X"00",X"55",X"A8",X"50",X"00",
		X"00",X"00",X"05",X"58",X"88",X"90",X"00",X"00",X"00",X"55",X"87",X"11",X"1E",X"00",X"00",X"05",
		X"58",X"71",X"17",X"75",X"00",X"00",X"05",X"58",X"89",X"77",X"59",X"00",X"00",X"09",X"58",X"88",
		X"55",X"59",X"A0",X"00",X"00",X"55",X"88",X"99",X"9F",X"A9",X"00",X"00",X"95",X"5F",X"FF",X"FA",
		X"95",X"00",X"00",X"05",X"55",X"59",X"99",X"59",X"00",X"00",X"09",X"55",X"55",X"99",X"9A",X"00",
		X"00",X"00",X"59",X"99",X"9A",X"90",X"00",X"00",X"00",X"95",X"99",X"A5",X"00",X"00",X"00",X"00",
		X"55",X"5A",X"50",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"99",X"55",X"59",X"00",X"00",
		X"9A",X"A5",X"55",X"00",X"00",X"A9",X"A0",X"55",X"00",X"00",X"A5",X"00",X"55",X"00",X"00",X"59",
		X"00",X"55",X"00",X"0A",X"5A",X"00",X"59",X"00",X"09",X"50",X"8A",X"50",X"00",X"05",X"55",X"89",
		X"50",X"00",X"89",X"58",X"85",X"5A",X"50",X"88",X"88",X"89",X"55",X"90",X"08",X"88",X"8A",X"50",
		X"00",X"00",X"08",X"88",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"99",X"55",X"55",
		X"90",X"00",X"00",X"9A",X"AA",X"55",X"55",X"00",X"00",X"A9",X"A0",X"00",X"55",X"A0",X"00",X"A5",
		X"00",X"09",X"59",X"00",X"00",X"95",X"00",X"09",X"50",X"00",X"00",X"59",X"00",X"A5",X"90",X"00",
		X"0A",X"50",X"00",X"A4",X"50",X"00",X"09",X"50",X"00",X"0A",X"45",X"00",X"05",X"55",X"90",X"00",
		X"A9",X"00",X"0A",X"58",X"88",X"00",X"00",X"00",X"08",X"88",X"88",X"88",X"80",X"00",X"00",X"88",
		X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"A9",X"55",X"50",X"00",X"00",X"00",
		X"00",X"00",X"A9",X"A0",X"A9",X"59",X"00",X"00",X"00",X"00",X"00",X"95",X"A0",X"0A",X"95",X"00",
		X"00",X"00",X"00",X"0A",X"55",X"00",X"00",X"55",X"00",X"00",X"00",X"D9",X"95",X"5A",X"00",X"00",
		X"55",X"0A",X"00",X"00",X"A4",X"50",X"00",X"00",X"00",X"95",X"95",X"00",X"00",X"04",X"50",X"00",
		X"00",X"00",X"A5",X"50",X"00",X"08",X"84",X"95",X"88",X"88",X"88",X"05",X"00",X"00",X"08",X"88",
		X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"55",X"55",X"50",X"00",X"00",X"99",X"55",X"59",X"00",X"00",X"9A",X"A5",X"55",X"00",X"00",
		X"AA",X"8A",X"55",X"00",X"0A",X"9A",X"A8",X"55",X"00",X"0A",X"49",X"A8",X"59",X"00",X"0A",X"45",
		X"09",X"5A",X"00",X"00",X"59",X"05",X"50",X"00",X"00",X"88",X"85",X"50",X"00",X"08",X"88",X"85",
		X"55",X"50",X"08",X"88",X"89",X"55",X"00",X"00",X"08",X"8A",X"50",X"00",X"55",X"55",X"50",X"00",
		X"00",X"99",X"55",X"55",X"A0",X"00",X"9A",X"A5",X"55",X"5A",X"00",X"A9",X"AA",X"A9",X"55",X"A0",
		X"0A",X"9A",X"8A",X"95",X"90",X"00",X"95",X"55",X"55",X"A0",X"00",X"54",X"59",X"00",X"00",X"00",
		X"54",X"50",X"00",X"00",X"0A",X"A9",X"50",X"00",X"00",X"09",X"AA",X"00",X"00",X"00",X"0A",X"95",
		X"A0",X"00",X"00",X"08",X"A5",X"58",X"80",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"88",X"88",
		X"88",X"00",X"00",X"00",X"88",X"80",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"09",X"55",X"55",
		X"50",X"00",X"00",X"09",X"99",X"55",X"55",X"90",X"00",X"0A",X"9A",X"A9",X"55",X"55",X"A0",X"00",
		X"AA",X"A0",X"0A",X"55",X"90",X"00",X"0A",X"9A",X"00",X"A5",X"90",X"00",X"00",X"A9",X"00",X"95",
		X"00",X"00",X"09",X"59",X"00",X"59",X"00",X"00",X"55",X"90",X"00",X"55",X"50",X"0A",X"5A",X"00",
		X"00",X"59",X"A0",X"00",X"39",X"88",X"80",X"00",X"00",X"00",X"A5",X"88",X"88",X"80",X"00",X"00",
		X"88",X"88",X"88",X"88",X"80",X"00",X"00",X"08",X"88",X"00",X"00",X"00",X"55",X"55",X"50",X"00",
		X"00",X"55",X"55",X"5A",X"00",X"00",X"99",X"55",X"5A",X"A0",X"00",X"0A",X"95",X"5A",X"A0",X"00",
		X"00",X"A5",X"5A",X"00",X"00",X"08",X"85",X"90",X"00",X"00",X"0A",X"55",X"A8",X"00",X"00",X"A5",
		X"58",X"88",X"00",X"0A",X"55",X"88",X"80",X"00",X"05",X"59",X"80",X"00",X"00",X"0A",X"95",X"50",
		X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"08",X"88",X"80",X"00",X"00",X"00",X"0E",X"11",X"17",
		X"00",X"00",X"00",X"00",X"05",X"77",X"11",X"70",X"FE",X"10",X"00",X"09",X"57",X"79",X"88",X"79",
		X"80",X"00",X"A9",X"55",X"58",X"88",X"95",X"00",X"09",X"AF",X"99",X"98",X"88",X"5A",X"00",X"05",
		X"9A",X"FF",X"FF",X"85",X"59",X"00",X"09",X"59",X"95",X"55",X"55",X"5A",X"00",X"0A",X"99",X"95",
		X"55",X"59",X"A0",X"00",X"00",X"9A",X"99",X"99",X"A0",X"00",X"00",X"00",X"05",X"A9",X"95",X"A0",
		X"00",X"00",X"00",X"00",X"5A",X"55",X"50",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"59",X"00",X"00",X"00",X"00",X"00",X"58",X"75",X"90",X"00",X"00",X"00",X"00",X"58",X"A5",
		X"50",X"00",X"00",X"00",X"00",X"98",X"88",X"55",X"00",X"00",X"00",X"0E",X"11",X"17",X"85",X"50",
		X"00",X"00",X"05",X"77",X"11",X"78",X"55",X"00",X"00",X"09",X"57",X"79",X"88",X"55",X"00",X"00",
		X"A9",X"55",X"58",X"88",X"59",X"00",X"09",X"AF",X"99",X"98",X"85",X"50",X"00",X"05",X"9A",X"FF",
		X"FF",X"55",X"90",X"00",X"09",X"59",X"99",X"55",X"55",X"00",X"00",X"0A",X"99",X"95",X"55",X"59",
		X"00",X"00",X"00",X"9A",X"99",X"99",X"50",X"00",X"00",X"00",X"05",X"A9",X"95",X"90",X"00",X"00",
		X"00",X"00",X"5A",X"55",X"50",X"00",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"02",
		X"66",X"66",X"62",X"00",X"00",X"00",X"06",X"63",X"66",X"66",X"00",X"00",X"00",X"06",X"60",X"06",
		X"63",X"00",X"00",X"00",X"06",X"60",X"06",X"60",X"00",X"00",X"00",X"05",X"60",X"06",X"60",X"00",
		X"00",X"00",X"00",X"66",X"05",X"63",X"00",X"00",X"00",X"00",X"66",X"00",X"66",X"00",X"00",X"00",
		X"06",X"66",X"00",X"66",X"00",X"00",X"00",X"66",X"38",X"88",X"66",X"88",X"00",X"08",X"88",X"88",
		X"36",X"66",X"88",X"80",X"00",X"88",X"88",X"66",X"38",X"88",X"00",X"00",X"08",X"88",X"88",X"88",
		X"80",X"00",X"00",X"00",X"88",X"88",X"88",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"03",
		X"86",X"66",X"60",X"00",X"00",X"03",X"66",X"63",X"00",X"00",X"00",X"02",X"66",X"00",X"00",X"00",
		X"00",X"06",X"60",X"00",X"00",X"00",X"00",X"05",X"62",X"00",X"00",X"00",X"00",X"03",X"26",X"60",
		X"00",X"00",X"00",X"00",X"32",X"63",X"88",X"80",X"00",X"06",X"28",X"66",X"88",X"88",X"00",X"66",
		X"33",X"63",X"88",X"80",X"00",X"00",X"06",X"68",X"88",X"00",X"00",X"00",X"00",X"88",X"00",X"00",
		X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"28",X"66",
		X"30",X"00",X"00",X"00",X"32",X"66",X"00",X"00",X"00",X"00",X"36",X"63",X"00",X"00",X"00",X"00",
		X"06",X"63",X"63",X"00",X"00",X"00",X"06",X"53",X"26",X"62",X"00",X"00",X"05",X"60",X"83",X"62",
		X"00",X"00",X"06",X"20",X"03",X"68",X"00",X"00",X"06",X"60",X"83",X"68",X"80",X"00",X"06",X"68",
		X"88",X"88",X"80",X"00",X"26",X"68",X"88",X"88",X"00",X"06",X"66",X"88",X"80",X"00",X"00",X"00",
		X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"06",X"66",X"66",X"62",X"00",X"00",X"00",X"66",X"63",
		X"66",X"66",X"00",X"00",X"06",X"62",X"00",X"06",X"63",X"00",X"00",X"25",X"60",X"00",X"06",X"60",
		X"00",X"00",X"36",X"66",X"20",X"09",X"60",X"00",X"00",X"00",X"36",X"60",X"03",X"66",X"00",X"00",
		X"00",X"06",X"20",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",X"66",X"00",X"00",X"08",X"88",
		X"88",X"36",X"66",X"80",X"00",X"00",X"08",X"88",X"66",X"38",X"88",X"00",X"00",X"00",X"08",X"88",
		X"88",X"80",X"00",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"00",X"06",X"66",X"66",
		X"62",X"00",X"00",X"00",X"00",X"66",X"63",X"66",X"66",X"00",X"00",X"00",X"02",X"66",X"00",X"26",
		X"63",X"00",X"00",X"00",X"05",X"60",X"00",X"06",X"60",X"00",X"00",X"00",X"06",X"20",X"00",X"06",
		X"63",X"23",X"00",X"00",X"06",X"20",X"00",X"05",X"62",X"26",X"00",X"00",X"06",X"60",X"00",X"00",
		X"00",X"66",X"00",X"00",X"06",X"60",X"00",X"00",X"00",X"63",X"00",X"03",X"66",X"68",X"88",X"88",
		X"88",X"88",X"00",X"06",X"63",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"88",X"88",X"88",X"00",
		X"00",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"06",X"86",X"66",X"60",X"00",X"00",
		X"00",X"36",X"36",X"66",X"00",X"00",X"00",X"00",X"63",X"66",X"68",X"00",X"00",X"00",X"00",X"53",
		X"66",X"33",X"60",X"00",X"00",X"00",X"00",X"66",X"32",X"68",X"00",X"00",X"00",X"00",X"66",X"86",
		X"88",X"80",X"00",X"00",X"00",X"56",X"60",X"88",X"88",X"80",X"00",X"00",X"00",X"66",X"00",X"88",
		X"88",X"00",X"00",X"00",X"06",X"68",X"88",X"80",X"00",X"00",X"00",X"36",X"28",X"88",X"80",X"00",
		X"00",X"00",X"66",X"88",X"88",X"80",X"00",X"00",X"66",X"66",X"60",X"00",X"06",X"86",X"66",X"60",
		X"00",X"02",X"66",X"66",X"00",X"00",X"26",X"66",X"00",X"00",X"00",X"56",X"33",X"26",X"30",X"00",
		X"66",X"66",X"66",X"60",X"00",X"02",X"30",X"06",X"60",X"00",X"06",X"68",X"83",X"60",X"00",X"06",
		X"68",X"88",X"00",X"00",X"36",X"68",X"88",X"88",X"00",X"66",X"38",X"88",X"88",X"80",X"08",X"88",
		X"88",X"88",X"00",X"00",X"00",X"03",X"61",X"11",X"63",X"00",X"00",X"00",X"00",X"06",X"76",X"66",
		X"66",X"00",X"00",X"00",X"00",X"06",X"88",X"88",X"66",X"00",X"00",X"00",X"00",X"06",X"86",X"88",
		X"63",X"30",X"00",X"00",X"00",X"03",X"82",X"88",X"86",X"60",X"00",X"00",X"00",X"63",X"88",X"85",
		X"36",X"66",X"00",X"00",X"02",X"35",X"71",X"66",X"23",X"26",X"30",X"00",X"03",X"77",X"86",X"66",
		X"66",X"66",X"60",X"03",X"57",X"E3",X"32",X"32",X"66",X"66",X"50",X"01",X"70",X"68",X"26",X"63",
		X"33",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"61",X"03",X"61",X"11",X"63",X"00",X"00",X"66",
		X"06",X"76",X"66",X"66",X"00",X"03",X"68",X"06",X"88",X"88",X"66",X"00",X"06",X"37",X"06",X"86",
		X"88",X"63",X"00",X"06",X"82",X"83",X"82",X"88",X"82",X"30",X"06",X"36",X"63",X"88",X"83",X"66",
		X"60",X"00",X"01",X"66",X"28",X"36",X"66",X"60",X"00",X"02",X"86",X"66",X"66",X"63",X"30",X"00",
		X"36",X"03",X"66",X"66",X"36",X"00",X"00",X"93",X"08",X"23",X"33",X"63",X"00",X"00",X"00",X"00",
		X"66",X"66",X"60",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"02",X"66",X"66",X"62",
		X"00",X"00",X"00",X"06",X"66",X"63",X"66",X"00",X"00",X"00",X"03",X"66",X"00",X"66",X"00",X"00",
		X"00",X"00",X"66",X"00",X"66",X"00",X"00",X"00",X"00",X"66",X"00",X"65",X"00",X"00",X"00",X"03",
		X"65",X"06",X"60",X"00",X"00",X"00",X"06",X"60",X"06",X"60",X"00",X"00",X"00",X"06",X"60",X"06",
		X"66",X"00",X"00",X"08",X"86",X"68",X"88",X"36",X"60",X"00",X"88",X"86",X"66",X"38",X"88",X"88",
		X"00",X"08",X"88",X"36",X"68",X"88",X"80",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",
		X"08",X"88",X"88",X"80",X"00",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"66",X"66",
		X"83",X"00",X"00",X"00",X"03",X"66",X"63",X"00",X"00",X"00",X"00",X"06",X"62",X"00",X"00",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"02",X"65",X"00",X"00",X"00",X"00",X"66",X"23",X"00",
		X"00",X"88",X"83",X"62",X"30",X"00",X"08",X"88",X"86",X"68",X"26",X"00",X"00",X"88",X"83",X"63",
		X"36",X"60",X"00",X"08",X"88",X"66",X"00",X"00",X"00",X"00",X"08",X"80",X"00",X"00",X"00",X"00",
		X"66",X"66",X"60",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"36",X"68",X"20",X"00",
		X"00",X"00",X"06",X"62",X"30",X"00",X"00",X"00",X"03",X"66",X"30",X"00",X"00",X"03",X"63",X"66",
		X"00",X"00",X"02",X"66",X"23",X"56",X"00",X"00",X"02",X"63",X"80",X"65",X"00",X"00",X"08",X"63",
		X"00",X"26",X"00",X"00",X"88",X"63",X"80",X"66",X"00",X"00",X"88",X"88",X"88",X"66",X"00",X"00",
		X"08",X"88",X"88",X"66",X"20",X"00",X"00",X"00",X"88",X"86",X"66",X"00",X"00",X"00",X"66",X"66",
		X"60",X"00",X"00",X"00",X"02",X"66",X"66",X"66",X"00",X"00",X"00",X"06",X"66",X"63",X"66",X"60",
		X"00",X"00",X"03",X"66",X"00",X"02",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"65",X"20",X"00",
		X"00",X"69",X"00",X"26",X"66",X"30",X"00",X"06",X"63",X"00",X"66",X"30",X"00",X"00",X"06",X"60",
		X"00",X"26",X"00",X"00",X"00",X"06",X"60",X"00",X"06",X"00",X"00",X"00",X"86",X"66",X"38",X"88",
		X"88",X"00",X"08",X"88",X"36",X"68",X"88",X"00",X"00",X"00",X"88",X"88",X"88",X"00",X"00",X"00",
		X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"00",X"02",X"66",X"66",X"66",X"00",X"00",X"00",
		X"00",X"06",X"66",X"63",X"66",X"60",X"00",X"00",X"00",X"03",X"66",X"20",X"06",X"62",X"00",X"00",
		X"00",X"00",X"66",X"00",X"00",X"65",X"00",X"00",X"03",X"23",X"66",X"00",X"00",X"26",X"00",X"00",
		X"06",X"22",X"65",X"00",X"00",X"26",X"00",X"00",X"06",X"60",X"00",X"00",X"00",X"66",X"00",X"00",
		X"03",X"60",X"00",X"00",X"00",X"66",X"00",X"00",X"08",X"88",X"88",X"88",X"88",X"66",X"63",X"00",
		X"00",X"08",X"88",X"88",X"88",X"83",X"66",X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"80",X"00",
		X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"00",X"66",X"66",X"86",X"00",X"00",X"00",
		X"00",X"06",X"66",X"36",X"30",X"00",X"00",X"00",X"08",X"66",X"63",X"60",X"00",X"00",X"00",X"63",
		X"36",X"63",X"50",X"00",X"00",X"08",X"62",X"36",X"60",X"00",X"00",X"00",X"88",X"86",X"86",X"60",
		X"00",X"00",X"88",X"88",X"80",X"66",X"50",X"00",X"08",X"88",X"80",X"06",X"60",X"00",X"00",X"00",
		X"88",X"88",X"66",X"00",X"00",X"00",X"00",X"88",X"88",X"26",X"30",X"00",X"00",X"00",X"88",X"88",
		X"86",X"60",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"66",X"66",X"86",X"00",X"00",X"06",
		X"66",X"62",X"00",X"00",X"00",X"06",X"66",X"20",X"00",X"36",X"23",X"36",X"50",X"00",X"66",X"66",
		X"66",X"60",X"00",X"66",X"00",X"32",X"00",X"00",X"63",X"88",X"66",X"00",X"00",X"08",X"88",X"66",
		X"00",X"08",X"88",X"88",X"66",X"30",X"88",X"88",X"88",X"36",X"60",X"08",X"88",X"88",X"88",X"00",
		X"00",X"03",X"61",X"11",X"63",X"00",X"00",X"00",X"00",X"06",X"66",X"66",X"76",X"00",X"00",X"00",
		X"00",X"06",X"68",X"88",X"86",X"00",X"00",X"00",X"00",X"33",X"68",X"86",X"86",X"00",X"00",X"00",
		X"00",X"66",X"88",X"82",X"83",X"00",X"00",X"00",X"06",X"66",X"35",X"88",X"83",X"60",X"00",X"00",
		X"36",X"23",X"26",X"61",X"75",X"32",X"00",X"00",X"66",X"66",X"66",X"66",X"87",X"73",X"00",X"00",
		X"56",X"66",X"62",X"32",X"33",X"E7",X"53",X"00",X"00",X"03",X"33",X"66",X"28",X"60",X"71",X"00",
		X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"03",X"61",X"11",X"63",X"01",X"60",X"00",X"06",X"66",X"66",X"76",X"06",
		X"60",X"00",X"06",X"68",X"88",X"86",X"08",X"63",X"00",X"03",X"68",X"86",X"86",X"07",X"36",X"00",
		X"32",X"88",X"82",X"83",X"82",X"86",X"00",X"66",X"63",X"88",X"83",X"66",X"36",X"00",X"66",X"66",
		X"38",X"26",X"61",X"00",X"00",X"33",X"66",X"66",X"66",X"82",X"00",X"00",X"06",X"36",X"66",X"63",
		X"06",X"30",X"00",X"03",X"63",X"33",X"28",X"03",X"90",X"00",X"00",X"66",X"66",X"60",X"00",X"00",
		X"00",X"00",X"66",X"66",X"60",X"00",X"02",X"66",X"66",X"20",X"00",X"06",X"66",X"33",X"20",X"00",
		X"06",X"60",X"36",X"30",X"00",X"06",X"60",X"06",X"30",X"00",X"06",X"60",X"05",X"60",X"00",X"05",
		X"60",X"03",X"63",X"00",X"00",X"63",X"80",X"62",X"00",X"00",X"66",X"86",X"66",X"00",X"63",X"66",
		X"88",X"62",X"80",X"36",X"66",X"88",X"88",X"80",X"00",X"63",X"88",X"88",X"00",X"00",X"08",X"88",
		X"00",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"26",X"66",X"66",X"20",X"00",X"06",X"66",
		X"66",X"33",X"20",X"00",X"26",X"60",X"00",X"36",X"30",X"00",X"05",X"62",X"00",X"06",X"30",X"00",
		X"00",X"62",X"00",X"06",X"20",X"00",X"00",X"66",X"30",X"05",X"60",X"00",X"00",X"64",X"30",X"00",
		X"63",X"00",X"06",X"43",X"00",X"00",X"66",X"00",X"03",X"30",X"00",X"36",X"66",X"00",X"00",X"00",
		X"08",X"88",X"63",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"08",X"88",X"88",X"80",X"00",
		X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"66",X"20",X"00",
		X"00",X"00",X"00",X"00",X"66",X"62",X"33",X"20",X"00",X"00",X"00",X"00",X"05",X"66",X"30",X"36",
		X"30",X"00",X"00",X"00",X"00",X"06",X"63",X"00",X"36",X"20",X"00",X"00",X"00",X"00",X"06",X"60",
		X"00",X"05",X"63",X"00",X"00",X"00",X"03",X"06",X"60",X"00",X"03",X"66",X"62",X"D0",X"00",X"06",
		X"66",X"20",X"00",X"00",X"00",X"64",X"30",X"00",X"00",X"66",X"30",X"00",X"00",X"00",X"64",X"00",
		X"00",X"00",X"06",X"08",X"88",X"88",X"86",X"24",X"88",X"00",X"00",X"00",X"08",X"88",X"88",X"88",
		X"88",X"88",X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"80",X"00",X"00",X"00",X"66",X"66",X"60",
		X"00",X"06",X"66",X"66",X"20",X"00",X"06",X"66",X"33",X"20",X"00",X"06",X"63",X"83",X"30",X"00",
		X"06",X"68",X"33",X"63",X"00",X"05",X"68",X"36",X"43",X"00",X"03",X"62",X"06",X"43",X"00",X"00",
		X"66",X"02",X"60",X"00",X"00",X"66",X"88",X"80",X"00",X"66",X"66",X"88",X"88",X"00",X"06",X"62",
		X"88",X"88",X"00",X"00",X"63",X"88",X"00",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"06",X"66",
		X"66",X"20",X"00",X"66",X"66",X"33",X"20",X"06",X"66",X"33",X"36",X"00",X"56",X"28",X"83",X"60",
		X"00",X"66",X"66",X"66",X"20",X"00",X"00",X"06",X"64",X"60",X"00",X"00",X"00",X"64",X"60",X"00",
		X"00",X"00",X"66",X"33",X"00",X"00",X"00",X"03",X"62",X"00",X"00",X"00",X"06",X"63",X"00",X"00",
		X"88",X"66",X"38",X"00",X"08",X"88",X"88",X"88",X"80",X"08",X"88",X"88",X"80",X"00",X"00",X"88",
		X"80",X"00",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"66",X"66",X"62",X"00",X"00",
		X"26",X"66",X"66",X"22",X"00",X"36",X"66",X"66",X"33",X"63",X"00",X"56",X"66",X"00",X"36",X"30",
		X"00",X"26",X"30",X"03",X"63",X"00",X"00",X"06",X"60",X"05",X"30",X"00",X"00",X"02",X"60",X"06",
		X"66",X"00",X"00",X"66",X"60",X"00",X"26",X"60",X"00",X"36",X"60",X"00",X"03",X"63",X"00",X"00",
		X"00",X"88",X"82",X"60",X"00",X"00",X"88",X"88",X"86",X"30",X"00",X"88",X"88",X"88",X"88",X"80",
		X"00",X"00",X"08",X"88",X"00",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"03",X"66",X"66",X"60",
		X"00",X"33",X"66",X"62",X"30",X"00",X"23",X"66",X"23",X"00",X"00",X"03",X"66",X"30",X"00",X"00",
		X"00",X"56",X"88",X"00",X"00",X"08",X"36",X"63",X"00",X"00",X"08",X"88",X"66",X"30",X"00",X"00",
		X"88",X"86",X"63",X"00",X"00",X"00",X"82",X"66",X"00",X"00",X"00",X"66",X"23",X"00",X"00",X"08",
		X"88",X"80",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"06",X"11",X"16",X"00",X"00",X"1E",
		X"00",X"61",X"17",X"76",X"60",X"00",X"87",X"58",X"88",X"76",X"66",X"60",X"00",X"08",X"71",X"88",
		X"66",X"66",X"20",X"00",X"00",X"87",X"A8",X"66",X"6F",X"26",X"00",X"00",X"06",X"5F",X"FF",X"F2",
		X"66",X"00",X"00",X"E6",X"86",X"66",X"63",X"66",X"00",X"00",X"68",X"66",X"66",X"62",X"6E",X"00",
		X"00",X"66",X"66",X"22",X"63",X"60",X"00",X"00",X"56",X"32",X"66",X"36",X"00",X"00",X"00",X"00",
		X"66",X"63",X"60",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",
		X"00",X"06",X"81",X"06",X"11",X"16",X"00",X"00",X"06",X"68",X"61",X"17",X"76",X"60",X"00",X"08",
		X"38",X"88",X"76",X"66",X"60",X"00",X"08",X"78",X"88",X"66",X"66",X"20",X"00",X"06",X"38",X"88",
		X"66",X"6F",X"26",X"00",X"06",X"66",X"8F",X"FF",X"F2",X"66",X"00",X"06",X"68",X"86",X"66",X"63",
		X"66",X"00",X"00",X"63",X"66",X"66",X"62",X"6E",X"00",X"00",X"66",X"66",X"22",X"63",X"60",X"00",
		X"00",X"56",X"32",X"66",X"36",X"00",X"00",X"00",X"00",X"66",X"63",X"60",X"00",X"00",X"00",X"66",
		X"66",X"60",X"00",X"00",X"26",X"66",X"62",X"00",X"00",X"23",X"36",X"66",X"00",X"00",X"36",X"30",
		X"66",X"00",X"00",X"36",X"00",X"66",X"00",X"00",X"65",X"00",X"66",X"00",X"03",X"63",X"00",X"65",
		X"00",X"02",X"60",X"83",X"60",X"00",X"06",X"66",X"86",X"60",X"00",X"82",X"68",X"86",X"63",X"60",
		X"88",X"88",X"86",X"66",X"30",X"08",X"88",X"83",X"60",X"00",X"00",X"08",X"88",X"00",X"00",X"00",
		X"66",X"66",X"60",X"00",X"00",X"00",X"26",X"66",X"66",X"20",X"00",X"00",X"23",X"36",X"66",X"66",
		X"00",X"00",X"36",X"30",X"00",X"66",X"20",X"00",X"36",X"00",X"02",X"65",X"00",X"00",X"26",X"00",
		X"02",X"60",X"00",X"00",X"65",X"00",X"36",X"60",X"00",X"03",X"60",X"00",X"34",X"60",X"00",X"06",
		X"60",X"00",X"03",X"46",X"00",X"06",X"66",X"30",X"00",X"33",X"00",X"03",X"68",X"88",X"00",X"00",
		X"00",X"08",X"88",X"88",X"88",X"80",X"00",X"00",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"26",X"66",X"66",X"00",X"00",X"00",X"00",
		X"00",X"00",X"23",X"32",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"36",X"30",X"36",X"65",X"00",
		X"00",X"00",X"00",X"00",X"26",X"30",X"03",X"66",X"00",X"00",X"00",X"00",X"03",X"65",X"00",X"00",
		X"66",X"00",X"00",X"00",X"D2",X"66",X"63",X"00",X"00",X"66",X"03",X"00",X"00",X"34",X"60",X"00",
		X"00",X"00",X"26",X"66",X"00",X"00",X"04",X"60",X"00",X"00",X"00",X"36",X"60",X"00",X"08",X"84",
		X"26",X"88",X"88",X"88",X"06",X"00",X"00",X"08",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"00",
		X"00",X"00",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"26",
		X"66",X"66",X"00",X"00",X"23",X"36",X"66",X"00",X"00",X"33",X"83",X"66",X"00",X"03",X"63",X"38",
		X"66",X"00",X"03",X"46",X"38",X"65",X"00",X"03",X"46",X"02",X"63",X"00",X"00",X"62",X"06",X"60",
		X"00",X"00",X"88",X"86",X"60",X"00",X"08",X"88",X"86",X"66",X"60",X"08",X"88",X"82",X"66",X"00",
		X"00",X"08",X"83",X"60",X"00",X"66",X"66",X"60",X"00",X"00",X"26",X"66",X"66",X"00",X"00",X"23",
		X"36",X"66",X"60",X"00",X"06",X"33",X"36",X"66",X"00",X"00",X"63",X"88",X"26",X"50",X"00",X"26",
		X"66",X"66",X"60",X"00",X"64",X"66",X"00",X"00",X"00",X"64",X"60",X"00",X"00",X"03",X"36",X"60",
		X"00",X"00",X"02",X"63",X"00",X"00",X"00",X"03",X"66",X"00",X"00",X"00",X"08",X"36",X"68",X"80",
		X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"88",X"88",X"88",X"00",X"00",X"00",X"88",X"80",X"00",
		X"00",X"66",X"66",X"60",X"00",X"00",X"02",X"66",X"66",X"60",X"00",X"00",X"02",X"26",X"66",X"66",
		X"20",X"00",X"03",X"63",X"36",X"66",X"66",X"30",X"00",X"36",X"30",X"06",X"66",X"50",X"00",X"03",
		X"63",X"00",X"36",X"20",X"00",X"00",X"35",X"00",X"66",X"00",X"00",X"06",X"66",X"00",X"62",X"00",
		X"00",X"66",X"20",X"00",X"66",X"60",X"03",X"63",X"00",X"00",X"66",X"30",X"00",X"62",X"88",X"80",
		X"00",X"00",X"00",X"36",X"88",X"88",X"80",X"00",X"00",X"88",X"88",X"88",X"88",X"80",X"00",X"00",
		X"08",X"88",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"66",X"66",X"63",X"00",X"00",X"32",
		X"66",X"63",X"30",X"00",X"03",X"26",X"63",X"20",X"00",X"00",X"36",X"63",X"00",X"00",X"08",X"86",
		X"50",X"00",X"00",X"03",X"66",X"38",X"00",X"00",X"36",X"68",X"88",X"00",X"03",X"66",X"88",X"80",
		X"00",X"06",X"62",X"80",X"00",X"00",X"03",X"26",X"60",X"00",X"00",X"00",X"88",X"88",X"00",X"00",
		X"08",X"88",X"80",X"00",X"00",X"00",X"06",X"11",X"16",X"00",X"00",X"00",X"00",X"66",X"77",X"11",
		X"60",X"0E",X"10",X"00",X"66",X"66",X"78",X"88",X"57",X"80",X"00",X"26",X"66",X"68",X"81",X"78",
		X"00",X"06",X"2F",X"66",X"68",X"A7",X"80",X"00",X"06",X"62",X"FF",X"FF",X"56",X"00",X"00",X"06",
		X"63",X"66",X"66",X"86",X"E0",X"00",X"0E",X"62",X"66",X"66",X"68",X"60",X"00",X"00",X"63",X"62",
		X"26",X"66",X"60",X"00",X"00",X"06",X"36",X"62",X"36",X"50",X"00",X"00",X"00",X"63",X"66",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"06",
		X"11",X"16",X"01",X"86",X"00",X"00",X"66",X"77",X"11",X"68",X"66",X"00",X"00",X"66",X"66",X"78",
		X"88",X"38",X"00",X"00",X"26",X"66",X"68",X"88",X"78",X"00",X"06",X"2F",X"66",X"68",X"88",X"36",
		X"00",X"06",X"62",X"FF",X"FF",X"86",X"66",X"00",X"06",X"63",X"66",X"66",X"88",X"66",X"00",X"0E",
		X"62",X"66",X"66",X"63",X"60",X"00",X"00",X"63",X"62",X"26",X"66",X"60",X"00",X"00",X"06",X"36",
		X"62",X"36",X"50",X"00",X"00",X"00",X"63",X"66",X"60",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"88",X"88",X"80",X"00",X"08",X"88",X"88",X"88",X"00",X"00",X"88",X"88",X"80",X"00",X"00",
		X"00",X"80",X"00",X"00",X"00",X"44",X"DD",X"CB",X"44",X"DD",X"CB",X"44",X"DD",X"00",X"00",X"0B",
		X"88",X"84",X"44",X"88",X"84",X"44",X"88",X"84",X"C0",X"00",X"C4",X"88",X"84",X"44",X"88",X"84",
		X"44",X"88",X"84",X"4B",X"00",X"44",X"88",X"84",X"44",X"88",X"84",X"44",X"88",X"84",X"44",X"00",
		X"44",X"88",X"84",X"44",X"88",X"84",X"44",X"88",X"84",X"44",X"00",X"44",X"44",X"DD",X"CB",X"44",
		X"DD",X"CB",X"44",X"DD",X"44",X"00",X"4B",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"C4",
		X"00",X"C8",X"47",X"24",X"88",X"88",X"88",X"88",X"47",X"24",X"8B",X"00",X"D8",X"24",X"4B",X"88",
		X"38",X"83",X"88",X"24",X"4B",X"84",X"00",X"48",X"B4",X"42",X"8E",X"E8",X"8E",X"E8",X"B4",X"42",
		X"84",X"00",X"48",X"42",X"74",X"8E",X"B8",X"8E",X"B8",X"42",X"74",X"8D",X"00",X"0B",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"C0",X"00",X"00",X"CD",X"44",X"BC",X"DD",X"44",X"BC",X"DD",
		X"4B",X"00",X"00",X"07",X"00",X"50",X"05",X"00",X"00",X"00",X"10",X"70",X"10",X"00",X"00",X"00",
		X"01",X"71",X"00",X"00",X"00",X"57",X"17",X"57",X"17",X"05",X"00",X"00",X"01",X"71",X"40",X"00",
		X"00",X"00",X"10",X"70",X"10",X"00",X"00",X"05",X"00",X"50",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"00",X"70",X"00",X"05",X"00",X"00",X"00",X"00",X"51",X"0A",X"19",X"A1",X"70",X"00",
		X"00",X"00",X"90",X"05",X"15",X"75",X"17",X"00",X"00",X"00",X"00",X"00",X"59",X"99",X"89",X"99",
		X"50",X"00",X"00",X"05",X"71",X"17",X"98",X"88",X"97",X"71",X"17",X"50",X"00",X"00",X"05",X"98",
		X"88",X"95",X"90",X"00",X"00",X"00",X"00",X"07",X"19",X"89",X"7A",X"00",X"90",X"00",X"00",X"00",
		X"71",X"A5",X"75",X"A1",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"10",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"90",X"70",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"09",X"99",X"00",X"97",X"00",X"00",
		X"00",X"00",X"00",X"90",X"00",X"99",X"99",X"8A",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"8A",X"88",X"A9",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"9A",X"A8",X"88",
		X"A8",X"90",X"00",X"00",X"00",X"00",X"05",X"71",X"59",X"88",X"88",X"88",X"88",X"A9",X"95",X"51",
		X"75",X"00",X"00",X"00",X"09",X"98",X"A8",X"88",X"8A",X"89",X"99",X"00",X"00",X"00",X"00",X"00",
		X"90",X"09",X"88",X"8A",X"88",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"9A",X"88",
		X"99",X"90",X"00",X"90",X"00",X"00",X"00",X"00",X"07",X"00",X"09",X"99",X"0A",X"59",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"48",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"8A",X"88",X"8A",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"8F",X"88",
		X"8A",X"89",X"00",X"00",X"00",X"00",X"08",X"A8",X"8A",X"88",X"88",X"88",X"88",X"88",X"80",X"00",
		X"00",X"00",X"08",X"88",X"88",X"8A",X"88",X"88",X"A8",X"F8",X"A8",X"A0",X"00",X"00",X"08",X"8A",
		X"8F",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"40",X"00",X"09",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"A8",X"F8",X"89",X"00",X"00",X"8A",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"80",X"00",X"08",X"8A",X"8F",X"8A",X"88",X"88",X"88",X"88",X"88",X"88",X"A0",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"8A",X"88",X"88",X"80",X"00",X"00",X"09",X"8A",X"88",X"8F",
		X"88",X"88",X"88",X"88",X"A8",X"80",X"00",X"00",X"00",X"08",X"8A",X"88",X"88",X"8F",X"88",X"8F",
		X"88",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A8",X"A8",X"84",X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"88",X"A8",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"80",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"50",X"07",X"00",X"00",X"00",X"10",X"70",X"10",X"00",X"00",X"00",
		X"01",X"71",X"00",X"00",X"05",X"07",X"17",X"57",X"17",X"50",X"00",X"00",X"41",X"71",X"00",X"00",
		X"00",X"00",X"10",X"70",X"10",X"00",X"00",X"05",X"00",X"50",X"05",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"05",X"00",X"00",X"00",X"05",
		X"00",X"00",X"70",X"00",X"70",X"00",X"00",X"00",X"00",X"71",X"A9",X"1A",X"01",X"50",X"00",X"00",
		X"00",X"00",X"07",X"15",X"75",X"15",X"00",X"90",X"00",X"00",X"00",X"59",X"99",X"89",X"99",X"50",
		X"00",X"00",X"57",X"11",X"77",X"98",X"88",X"97",X"11",X"75",X"00",X"00",X"00",X"95",X"98",X"88",
		X"95",X"00",X"00",X"00",X"00",X"90",X"0A",X"79",X"89",X"17",X"00",X"00",X"00",X"00",X"00",X"01",
		X"A5",X"75",X"A1",X"70",X"00",X"00",X"00",X"00",X"10",X"00",X"10",X"00",X"05",X"00",X"00",X"00",
		X"05",X"00",X"00",X"70",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"90",X"09",X"99",X"09",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"9A",X"89",X"99",X"90",X"00",X"90",X"00",X"00",X"00",X"00",
		X"90",X"99",X"A8",X"8A",X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"A8",X"88",
		X"AA",X"99",X"00",X"00",X"00",X"05",X"71",X"55",X"99",X"A8",X"88",X"88",X"88",X"89",X"51",X"75",
		X"00",X"00",X"00",X"09",X"99",X"8A",X"88",X"88",X"A8",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"98",X"8A",X"88",X"89",X"00",X"90",X"00",X"00",X"00",X"00",X"90",X"00",X"99",X"98",X"8A",
		X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"5A",X"09",X"99",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"8A",X"88",X"8A",X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"8A",X"88",X"8F",
		X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"8A",X"88",X"A8",
		X"00",X"00",X"00",X"A8",X"A8",X"F8",X"A8",X"88",X"8A",X"88",X"88",X"88",X"00",X"00",X"48",X"88",
		X"88",X"88",X"88",X"88",X"88",X"8F",X"8A",X"88",X"00",X"09",X"88",X"F8",X"A8",X"88",X"88",X"88",
		X"88",X"88",X"88",X"89",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"8A",X"80",
		X"00",X"A8",X"88",X"88",X"88",X"88",X"88",X"8A",X"8F",X"8A",X"88",X"00",X"00",X"88",X"88",X"8A",
		X"88",X"88",X"88",X"88",X"88",X"88",X"80",X"00",X"00",X"88",X"A8",X"88",X"88",X"88",X"8F",X"88",
		X"8A",X"89",X"00",X"00",X"00",X"08",X"8F",X"88",X"8F",X"88",X"88",X"8A",X"88",X"00",X"00",X"00",
		X"00",X"00",X"08",X"88",X"88",X"88",X"88",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"84",X"88",X"A8",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"A8",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"DC",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"4D",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"44",X"48",X"88",X"84",
		X"00",X"00",X"00",X"00",X"00",X"00",X"8C",X"CB",X"D8",X"88",X"88",X"88",X"DC",X"00",X"00",X"00",
		X"00",X"08",X"47",X"24",X"44",X"88",X"88",X"44",X"4D",X"B0",X"00",X"00",X"00",X"08",X"24",X"4B",
		X"88",X"48",X"44",X"44",X"48",X"84",X"40",X"00",X"00",X"08",X"B4",X"42",X"88",X"DC",X"44",X"48",
		X"88",X"88",X"8D",X"C0",X"00",X"08",X"42",X"74",X"88",X"8D",X"B4",X"88",X"88",X"88",X"44",X"DB",
		X"00",X"00",X"BD",X"88",X"EE",X"38",X"88",X"44",X"88",X"44",X"44",X"48",X"40",X"00",X"0C",X"D8",
		X"EB",X"88",X"38",X"88",X"DC",X"44",X"48",X"88",X"40",X"00",X"00",X"88",X"88",X"8E",X"E8",X"88",
		X"8D",X"B8",X"88",X"88",X"40",X"00",X"00",X"08",X"88",X"8E",X"B8",X"47",X"24",X"88",X"88",X"88",
		X"C0",X"00",X"00",X"00",X"08",X"88",X"88",X"24",X"4B",X"88",X"88",X"4C",X"00",X"00",X"00",X"00",
		X"00",X"8B",X"D8",X"B4",X"42",X"88",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"42",
		X"74",X"8B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"48",X"84",X"DC",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"84",X"44",X"44",X"84",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"8D",X"C4",X"44",X"88",X"88",X"84",X"00",X"00",X"00",X"00",X"08",X"42",X"74",
		X"DB",X"88",X"88",X"88",X"8D",X"C0",X"00",X"00",X"00",X"0D",X"B4",X"42",X"88",X"48",X"88",X"84",
		X"44",X"DB",X"40",X"00",X"00",X"0B",X"24",X"4B",X"88",X"84",X"84",X"44",X"44",X"88",X"84",X"00",
		X"00",X"0C",X"47",X"24",X"88",X"88",X"DC",X"44",X"88",X"88",X"88",X"DC",X"00",X"00",X"D8",X"88",
		X"EE",X"38",X"8D",X"B4",X"88",X"88",X"84",X"4D",X"B0",X"00",X"08",X"88",X"BE",X"88",X"38",X"88",
		X"48",X"84",X"44",X"44",X"40",X"00",X"00",X"88",X"88",X"8E",X"E8",X"88",X"8D",X"C4",X"44",X"88",
		X"40",X"00",X"00",X"08",X"88",X"8B",X"E8",X"42",X"74",X"DB",X"88",X"88",X"40",X"00",X"00",X"00",
		X"0B",X"D8",X"88",X"B4",X"42",X"88",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"CD",X"88",X"24",
		X"4B",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"47",X"24",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"8B",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"C0",X"00",X"00",X"00",X"00",X"20",X"49",X"4E",X"46",X"45",X"52",X"4E",
		X"4F",X"20",X"2D",X"20",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"28",X"43",
		X"29",X"20",X"31",X"39",X"38",X"34",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",
		X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",
		X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",
		X"88",X"8D",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"88",X"88",X"44",X"DB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"48",X"44",X"44",X"48",X"44",X"00",X"00",X"00",X"00",
		X"0D",X"4B",X"24",X"DC",X"44",X"48",X"88",X"88",X"D0",X"00",X"00",X"00",X"0B",X"24",X"47",X"8D",
		X"B8",X"88",X"88",X"88",X"4C",X"D0",X"00",X"00",X"0C",X"74",X"42",X"88",X"88",X"48",X"88",X"44",
		X"44",X"B4",X"00",X"00",X"0D",X"42",X"B4",X"88",X"88",X"8D",X"C4",X"44",X"48",X"88",X"48",X"00",
		X"00",X"88",X"88",X"BE",X"38",X"88",X"DB",X"48",X"88",X"88",X"8C",X"D0",X"00",X"08",X"88",X"EE",
		X"88",X"38",X"88",X"84",X"88",X"88",X"44",X"B0",X"00",X"00",X"8D",X"88",X"8B",X"E8",X"88",X"88",
		X"D8",X"44",X"44",X"D0",X"00",X"00",X"0B",X"C8",X"8E",X"E8",X"4B",X"24",X"8C",X"44",X"48",X"40",
		X"00",X"00",X"00",X"0D",X"88",X"88",X"24",X"47",X"8B",X"48",X"88",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"74",X"42",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"42",X"B4",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"C0",X"88",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BD",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"88",X"84",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"88",X"88",X"88",X"DC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"BC",X"88",X"48",X"88",X"84",X"4D",X"BD",X"00",X"00",X"00",X"00",X"0C",X"42",X"B4",X"84",
		X"84",X"44",X"44",X"88",X"40",X"00",X"00",X"00",X"0D",X"74",X"42",X"8D",X"E4",X"44",X"88",X"88",
		X"8D",X"D0",X"00",X"00",X"08",X"24",X"47",X"88",X"DB",X"48",X"88",X"88",X"84",X"CB",X"00",X"00",
		X"08",X"4B",X"24",X"88",X"88",X"84",X"88",X"84",X"44",X"44",X"84",X"00",X"00",X"88",X"88",X"EB",
		X"38",X"88",X"DC",X"44",X"44",X"88",X"88",X"40",X"00",X"0C",X"D8",X"EE",X"88",X"38",X"8D",X"B4",
		X"88",X"88",X"88",X"C0",X"00",X"00",X"BD",X"88",X"8E",X"B8",X"88",X"88",X"48",X"88",X"84",X"B0",
		X"00",X"00",X"08",X"88",X"8E",X"E8",X"42",X"B4",X"84",X"84",X"4D",X"40",X"00",X"00",X"00",X"08",
		X"88",X"88",X"74",X"42",X"8D",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"24",X"47",
		X"8B",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"4B",X"24",X"8C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"D8",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"44",X"44",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"44",X"44",
		X"40",X"00",X"00",X"00",X"00",X"04",X"44",X"08",X"44",X"44",X"44",X"80",X"00",X"00",X"00",X"04",
		X"40",X"00",X"44",X"84",X"44",X"48",X"40",X"00",X"00",X"00",X"04",X"48",X"88",X"84",X"48",X"88",
		X"84",X"40",X"00",X"00",X"00",X"00",X"48",X"80",X"84",X"44",X"44",X"44",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"44",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"84",
		X"44",X"40",X"40",X"00",X"44",X"40",X"00",X"00",X"00",X"08",X"88",X"88",X"80",X"04",X"04",X"44",
		X"40",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"84",X"44",X"84",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"84",X"44",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"44",X"48",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"BC",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4D",X"44",
		X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"88",X"88",X"44",X"44",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"D8",X"88",X"88",X"88",X"DB",X"CC",X"80",X"00",X"00",X"00",X"00",
		X"BD",X"44",X"48",X"88",X"84",X"44",X"27",X"48",X"00",X"00",X"00",X"44",X"88",X"44",X"44",X"48",
		X"48",X"8B",X"44",X"28",X"00",X"00",X"CD",X"88",X"88",X"88",X"44",X"4C",X"D8",X"82",X"44",X"B8",
		X"00",X"0B",X"D4",X"48",X"88",X"88",X"84",X"BD",X"88",X"84",X"72",X"48",X"00",X"48",X"44",X"44",
		X"48",X"84",X"48",X"88",X"3E",X"E8",X"8D",X"B0",X"00",X"48",X"88",X"44",X"4C",X"D8",X"88",X"38",
		X"8B",X"E8",X"DC",X"00",X"00",X"48",X"88",X"88",X"BD",X"88",X"88",X"EE",X"88",X"88",X"80",X"00",
		X"00",X"C8",X"88",X"88",X"84",X"27",X"48",X"BE",X"88",X"88",X"00",X"00",X"00",X"0C",X"48",X"88",
		X"8B",X"44",X"28",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"D8",X"82",X"44",X"B8",X"DB",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"84",X"72",X"4D",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C8",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BC",X"D4",X"88",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"84",X"44",X"44",X"88",X"80",X"00",X"00",X"00",X"00",X"00",
		X"04",X"88",X"88",X"84",X"44",X"CD",X"88",X"80",X"00",X"00",X"00",X"00",X"CD",X"88",X"88",X"88",
		X"8B",X"D4",X"72",X"48",X"00",X"00",X"00",X"4B",X"D4",X"44",X"88",X"88",X"48",X"82",X"44",X"BD",
		X"00",X"00",X"04",X"88",X"84",X"44",X"44",X"84",X"88",X"8B",X"44",X"2B",X"00",X"0C",X"D8",X"88",
		X"88",X"84",X"4C",X"D8",X"88",X"84",X"27",X"4C",X"00",X"BD",X"44",X"88",X"88",X"84",X"BD",X"88",
		X"3E",X"E8",X"88",X"D0",X"00",X"44",X"44",X"44",X"88",X"48",X"88",X"38",X"8E",X"B8",X"88",X"00",
		X"00",X"48",X"84",X"44",X"CD",X"88",X"88",X"EE",X"88",X"88",X"80",X"00",X"00",X"48",X"88",X"8B",
		X"D4",X"72",X"48",X"EB",X"88",X"88",X"00",X"00",X"00",X"00",X"88",X"88",X"82",X"44",X"B8",X"88",
		X"DB",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"8B",X"44",X"28",X"8D",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"84",X"27",X"48",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DB",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"88",X"84",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"D4",X"48",X"88",X"84",X"40",X"00",X"00",X"00",X"00",X"00",X"04",X"48",X"44",X"44",
		X"48",X"48",X"88",X"80",X"00",X"00",X"00",X"00",X"D8",X"88",X"88",X"44",X"4C",X"D4",X"2B",X"4D",
		X"00",X"00",X"00",X"DC",X"48",X"88",X"88",X"88",X"BD",X"87",X"44",X"2B",X"00",X"00",X"04",X"B4",
		X"44",X"48",X"88",X"48",X"88",X"82",X"44",X"7C",X"00",X"08",X"48",X"88",X"44",X"44",X"CD",X"88",
		X"88",X"84",X"B2",X"4D",X"00",X"DC",X"88",X"88",X"88",X"4B",X"D8",X"88",X"3E",X"B8",X"88",X"80",
		X"00",X"B4",X"48",X"88",X"84",X"88",X"88",X"38",X"8E",X"E8",X"88",X"00",X"00",X"D4",X"44",X"48",
		X"D8",X"88",X"88",X"EB",X"88",X"8D",X"80",X"00",X"00",X"48",X"44",X"4C",X"84",X"2B",X"48",X"EE",
		X"88",X"CB",X"00",X"00",X"00",X"08",X"88",X"4B",X"87",X"44",X"28",X"88",X"8D",X"00",X"00",X"00",
		X"00",X"00",X"08",X"88",X"82",X"44",X"78",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"84",X"B2",X"48",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"80",X"C8",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DB",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4D",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"84",X"88",X"84",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"D8",X"88",
		X"88",X"84",X"40",X"00",X"00",X"00",X"00",X"00",X"0D",X"BD",X"44",X"88",X"88",X"48",X"8C",X"B0",
		X"00",X"00",X"00",X"00",X"48",X"84",X"44",X"44",X"84",X"84",X"B2",X"4C",X"00",X"00",X"00",X"DD",
		X"88",X"88",X"84",X"44",X"ED",X"82",X"44",X"7D",X"00",X"00",X"0B",X"C4",X"88",X"88",X"88",X"4B",
		X"D8",X"87",X"44",X"28",X"00",X"04",X"84",X"44",X"44",X"88",X"84",X"88",X"88",X"84",X"2B",X"48",
		X"00",X"48",X"88",X"84",X"44",X"4C",X"D8",X"88",X"3B",X"E8",X"88",X"80",X"00",X"C8",X"88",X"88",
		X"84",X"BD",X"88",X"38",X"8E",X"E8",X"DC",X"00",X"00",X"B4",X"88",X"88",X"48",X"88",X"88",X"BE",
		X"88",X"8D",X"B0",X"00",X"00",X"4D",X"44",X"84",X"84",X"B2",X"48",X"EE",X"88",X"88",X"00",X"00",
		X"00",X"04",X"44",X"4D",X"82",X"44",X"78",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"04",X"4B",
		X"87",X"44",X"28",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"84",X"2B",X"4D",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"DB",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"44",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"44",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"44",X"44",X"48",
		X"04",X"44",X"00",X"00",X"00",X"00",X"00",X"48",X"44",X"44",X"84",X"40",X"00",X"44",X"00",X"00",
		X"00",X"00",X"44",X"88",X"88",X"44",X"88",X"88",X"44",X"00",X"00",X"00",X"00",X"44",X"44",X"44",
		X"44",X"80",X"88",X"40",X"00",X"00",X"00",X"00",X"04",X"44",X"44",X"48",X"80",X"00",X"00",X"00",
		X"44",X"40",X"00",X"40",X"44",X"44",X"88",X"80",X"00",X"00",X"00",X"44",X"44",X"04",X"00",X"88",
		X"88",X"88",X"00",X"00",X"00",X"00",X"04",X"84",X"44",X"88",X"88",X"88",X"80",X"00",X"00",X"00",
		X"00",X"00",X"08",X"84",X"44",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"44",
		X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"B4",X"44",X"44",X"44",X"44",X"B0",X"C4",X"44",X"44",X"44",X"44",X"C0",X"D4",X"44",
		X"44",X"44",X"44",X"D0",X"D8",X"88",X"88",X"88",X"88",X"D0",X"48",X"88",X"88",X"88",X"88",X"40",
		X"48",X"88",X"88",X"88",X"88",X"40",X"B4",X"44",X"44",X"44",X"44",X"B0",X"C4",X"44",X"44",X"44",
		X"44",X"C0",X"D4",X"44",X"44",X"44",X"44",X"D0",X"D8",X"88",X"88",X"88",X"88",X"D0",X"48",X"88",
		X"88",X"88",X"88",X"40",X"48",X"88",X"88",X"88",X"88",X"40",X"B4",X"44",X"44",X"44",X"44",X"B0",
		X"C4",X"44",X"44",X"44",X"44",X"C0",X"D4",X"44",X"44",X"44",X"44",X"D0",X"D8",X"88",X"88",X"88",
		X"88",X"D0",X"48",X"88",X"88",X"88",X"88",X"40",X"48",X"88",X"88",X"88",X"88",X"40",X"B4",X"44",
		X"44",X"44",X"44",X"B0",X"00",X"BB",X"B0",X"00",X"0C",X"B1",X"BC",X"00",X"00",X"BB",X"B0",X"00",
		X"00",X"11",X"10",X"00",X"01",X"11",X"11",X"00",X"00",X"11",X"10",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CB",X"C4",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"CB",X"8B",X"BB",X"CD",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",
		X"48",X"88",X"8C",X"CB",X"BB",X"CD",X"00",X"0B",X"00",X"00",X"00",X"04",X"5F",X"88",X"88",X"8B",
		X"C4",X"D0",X"DB",X"00",X"00",X"00",X"0D",X"32",X"24",X"5F",X"88",X"47",X"BB",X"BC",X"00",X"00",
		X"00",X"02",X"23",X"44",X"88",X"8C",X"4C",X"BC",X"CD",X"00",X"00",X"03",X"22",X"44",X"44",X"BC",
		X"CB",X"4D",X"CC",X"D0",X"00",X"04",X"36",X"34",X"48",X"AB",X"7B",X"BC",X"D4",X"00",X"00",X"00",
		X"36",X"24",X"48",X"88",X"88",X"BB",X"CD",X"DD",X"00",X"00",X"00",X"38",X"34",X"80",X"CC",X"C8",
		X"8B",X"DD",X"D0",X"00",X"00",X"00",X"43",X"40",X"00",X"BB",X"BB",X"8D",X"DD",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"BB",X"BD",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CB",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"91",X"60",X"00",X"00",X"A9",X"11",X"1A",
		X"00",X"00",X"97",X"57",X"90",X"00",X"09",X"A0",X"A0",X"00",X"00",X"00",X"90",X"00",X"5A",X"00",
		X"60",X"00",X"00",X"07",X"E9",X"18",X"65",X"A0",X"00",X"0A",X"09",X"A8",X"88",X"89",X"57",X"00",
		X"0E",X"5A",X"81",X"88",X"15",X"00",X"00",X"A0",X"98",X"9F",X"97",X"00",X"70",X"00",X"00",X"E5",
		X"09",X"00",X"90",X"00",X"00",X"0A",X"0A",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"00",X"00",X"00",X"00",X"A0",X"05",X"00",X"00",X"60",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"50",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"09",X"00",X"50",X"90",X"0E",X"00",X"A0",X"0E",X"00",X"A0",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"B0",X"00",X"00",
		X"0B",X"00",X"00",X"00",X"00",X"00",X"04",X"CB",X"C0",X"00",X"00",X"0B",X"00",X"00",X"00",X"0D",
		X"CB",X"BB",X"8B",X"C0",X"00",X"00",X"0B",X"00",X"0D",X"CB",X"BB",X"CC",X"88",X"88",X"40",X"00",
		X"00",X"0B",X"D0",X"D4",X"CB",X"88",X"88",X"8F",X"54",X"00",X"00",X"00",X"0C",X"BB",X"B7",X"48",
		X"8F",X"54",X"22",X"3D",X"00",X"00",X"00",X"0D",X"CC",X"BC",X"4C",X"88",X"84",X"43",X"22",X"00",
		X"00",X"00",X"00",X"DC",X"CD",X"4B",X"CC",X"B4",X"44",X"42",X"23",X"00",X"00",X"00",X"00",X"04",
		X"DC",X"BB",X"7B",X"A8",X"44",X"36",X"34",X"00",X"00",X"00",X"0D",X"DD",X"CB",X"B8",X"88",X"88",
		X"44",X"26",X"30",X"00",X"00",X"00",X"DD",X"DB",X"88",X"CC",X"C0",X"84",X"38",X"30",X"00",X"00",
		X"00",X"0D",X"DD",X"8B",X"BB",X"B0",X"00",X"43",X"40",X"00",X"00",X"00",X"00",X"DD",X"BB",X"BC",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DB",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"61",X"99",X"00",X"00",X"0A",X"11",X"19",X"A0",X"00",X"00",X"97",X"57",X"90",X"00",X"00",X"00",
		X"A0",X"A9",X"00",X"00",X"60",X"0A",X"50",X"00",X"90",X"00",X"00",X"A5",X"68",X"19",X"E7",X"00",
		X"00",X"07",X"59",X"88",X"88",X"A9",X"0A",X"00",X"00",X"05",X"18",X"81",X"8A",X"5E",X"00",X"00",
		X"70",X"07",X"9F",X"98",X"90",X"A0",X"00",X"00",X"90",X"09",X"05",X"E0",X"00",X"00",X"00",X"00",
		X"50",X"0A",X"0A",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"05",
		X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"A0",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"90",X"50",X"09",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"A0",X"0E",
		X"00",X"A0",X"0E",X"00",X"00",X"00",X"00",X"F0",X"00",X"0F",X"00",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"0B",X"BB",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"B0",X"B0",X"00",X"90",X"00",X"00",X"0C",X"0B",X"BC",X"00",X"00",X"00",X"B0",
		X"CB",X"D0",X"00",X"07",X"00",X"C0",X"00",X"00",X"D0",X"00",X"00",X"B0",X"0B",X"00",X"00",X"00",
		X"10",X"70",X"10",X"70",X"0D",X"00",X"DC",X"B0",X"00",X"05",X"00",X"00",X"01",X"11",X"00",X"00",
		X"00",X"0C",X"CB",X"00",X"02",X"00",X"00",X"51",X"11",X"81",X"11",X"79",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"C0",X"00",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"07",X"00",
		X"10",X"70",X"10",X"09",X"00",X"C0",X"00",X"00",X"02",X"40",X"0D",X"00",X"00",X"C0",X"07",X"00",
		X"0D",X"00",X"00",X"00",X"00",X"00",X"23",X"00",X"0B",X"00",X"00",X"0D",X"DD",X"00",X"00",X"00",
		X"04",X"02",X"34",X"0C",X"00",X"0B",X"CC",X"00",X"DD",X"00",X"00",X"00",X"00",X"06",X"30",X"00",
		X"00",X"00",X"B0",X"0D",X"D0",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"BB",X"BD",X"00",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"D0",X"0D",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"79",X"00",
		X"70",X"09",X"10",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"01",X"99",X"19",X"91",
		X"00",X"70",X"00",X"00",X"00",X"D0",X"0D",X"00",X"00",X"00",X"09",X"99",X"89",X"99",X"00",X"00",
		X"00",X"00",X"00",X"D0",X"00",X"05",X"00",X"00",X"91",X"98",X"88",X"91",X"90",X"00",X"00",X"00",
		X"00",X"D0",X"00",X"00",X"05",X"11",X"19",X"88",X"88",X"89",X"11",X"17",X"90",X"00",X"0D",X"00",
		X"30",X"00",X"00",X"00",X"91",X"98",X"88",X"91",X"90",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"00",X"00",X"09",X"99",X"89",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"07",X"00",
		X"01",X"99",X"19",X"91",X"00",X"09",X"00",X"D0",X"00",X"00",X"03",X"00",X"00",X"00",X"19",X"00",
		X"70",X"09",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"0B",X"00",X"00",X"D0",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"03",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"0A",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",
		X"00",X"70",X"A0",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"A0",X"09",X"89",X"00",
		X"01",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"0A",X"99",X"98",X"88",X"99",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"88",X"89",X"88",X"90",X"0A",X"00",X"00",X"00",X"00",
		X"0A",X"A0",X"0A",X"99",X"88",X"88",X"89",X"90",X"00",X"00",X"A0",X"00",X"90",X"00",X"00",X"A9",
		X"88",X"88",X"88",X"88",X"89",X"A0",X"00",X"00",X"00",X"00",X"97",X"19",X"98",X"88",X"88",X"88",
		X"88",X"88",X"99",X"17",X"A0",X"00",X"00",X"00",X"0A",X"A9",X"89",X"88",X"88",X"89",X"89",X"AA",
		X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"98",X"88",X"88",X"88",X"90",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"0A",X"98",X"A8",X"89",X"88",X"90",X"09",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"0A",X"99",X"98",X"88",X"99",X"9A",X"00",X"0A",X"00",X"00",X"00",X"05",X"00",X"01",X"00",X"09",
		X"89",X"00",X"0A",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"0A",X"0A",X"90",X"0A",X"00",
		X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"A0",X"09",X"00",X"A0",
		X"00",X"90",X"00",X"E0",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"A0",X"00",X"00",X"00",X"00",X"0F",X"00",X"A0",X"00",X"A0",X"00",X"00",X"A0",X"00",X"F0",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"00",X"0E",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"09",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"A0",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"0A",X"00",
		X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"A0",X"0A",X"00",
		X"00",X"A0",X"00",X"A0",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"B0",X"00",X"00",X"00",X"00",X"00",X"CB",X"BB",X"00",X"00",X"00",X"B0",
		X"B0",X"00",X"00",X"0C",X"BB",X"0C",X"00",X"00",X"00",X"90",X"00",X"B0",X"B0",X"00",X"00",X"D0",
		X"00",X"00",X"C0",X"07",X"00",X"00",X"DB",X"C0",X"BC",X"D0",X"0D",X"00",X"70",X"10",X"70",X"10",
		X"00",X"00",X"0B",X"00",X"0B",X"CC",X"00",X"00",X"00",X"01",X"11",X"00",X"00",X"05",X"00",X"00",
		X"00",X"B0",X"00",X"09",X"71",X"11",X"81",X"11",X"50",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"11",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"C0",X"09",X"00",X"10",X"70",X"10",
		X"07",X"00",X"20",X"00",X"00",X"00",X"0D",X"00",X"07",X"00",X"C0",X"00",X"0D",X"00",X"42",X"00",
		X"00",X"00",X"0D",X"DD",X"00",X"00",X"0B",X"00",X"03",X"20",X"00",X"00",X"00",X"00",X"0D",X"D0",
		X"0C",X"CB",X"00",X"0C",X"04",X"32",X"04",X"00",X"00",X"00",X"00",X"DD",X"00",X"B0",X"00",X"00",
		X"00",X"36",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"0D",X"BB",X"BC",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"DB",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"00",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"70",X"09",X"70",
		X"00",X"00",X"00",X"D0",X"D0",X"00",X"00",X"00",X"70",X"01",X"99",X"19",X"91",X"00",X"00",X"00",
		X"00",X"D0",X"D0",X"00",X"00",X"00",X"00",X"09",X"99",X"89",X"99",X"00",X"00",X"00",X"0D",X"00",
		X"D0",X"00",X"00",X"00",X"00",X"91",X"98",X"88",X"91",X"90",X"00",X"05",X"00",X"00",X"0D",X"00",
		X"00",X"97",X"11",X"19",X"88",X"88",X"89",X"11",X"15",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",
		X"00",X"91",X"98",X"88",X"91",X"90",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"09",
		X"99",X"89",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"09",X"00",X"01",X"99",X"19",
		X"91",X"00",X"07",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"00",X"70",X"09",X"10",
		X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"D0",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"D0",X"00",X"0B",X"00",X"00",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"0A",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"A0",X"70",X"00",X"00",
		X"50",X"00",X"00",X"00",X"00",X"00",X"50",X"01",X"00",X"09",X"89",X"00",X"A1",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"98",X"88",X"99",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"00",X"98",X"89",X"88",X"88",X"90",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"99",
		X"88",X"88",X"89",X"9A",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"A9",X"88",X"88",X"88",X"88",
		X"89",X"A0",X"00",X"00",X"90",X"00",X"A7",X"19",X"98",X"88",X"88",X"88",X"88",X"88",X"99",X"17",
		X"90",X"00",X"00",X"00",X"0A",X"A9",X"89",X"88",X"88",X"89",X"89",X"AA",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"98",X"88",X"88",X"88",X"90",X"00",X"00",X"0A",X"00",X"00",X"00",X"09",X"00",
		X"98",X"89",X"88",X"A8",X"9A",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"0A",X"99",X"98",X"88",
		X"99",X"9A",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"1A",X"00",X"09",X"89",X"00",X"01",X"00",
		X"05",X"00",X"00",X"00",X"00",X"05",X"00",X"0A",X"00",X"9A",X"0A",X"00",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"A0",X"00",X"E0",X"00",X"90",X"00",X"A0",
		X"09",X"00",X"A0",X"00",X"00",X"00",X"00",X"A0",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"F0",X"00",X"A0",X"00",X"00",X"A0",X"00",X"A0",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"0E",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"A9",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"09",X"A0",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"0F",X"00",
		X"0A",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"A0",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"09",X"00",X"0A",X"00",X"00",X"A0",X"00",X"00",X"A0",X"00",X"A0",X"00",X"0A",
		X"00",X"A0",X"00",X"00",X"06",X"00",X"0E",X"00",X"0F",X"00",X"01",X"00",X"06",X"00",X"0E",X"00",
		X"0F",X"00",X"01",X"00",X"0E",X"00",X"0F",X"00",X"01",X"00",X"06",X"00",X"0E",X"00",X"0F",X"00",
		X"01",X"00",X"06",X"00",X"0F",X"00",X"01",X"00",X"06",X"00",X"0E",X"00",X"0F",X"00",X"01",X"00",
		X"06",X"00",X"0E",X"00",X"01",X"00",X"06",X"00",X"0E",X"00",X"0F",X"00",X"01",X"00",X"06",X"00",
		X"0E",X"00",X"0F",X"00",X"36",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"32",X"46",
		X"30",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"32",X"22",X"40",X"00",X"00",X"00",X"00",
		X"B0",X"00",X"00",X"04",X"32",X"23",X"00",X"00",X"00",X"0D",X"BC",X"00",X"00",X"00",X"43",X"32",
		X"28",X"CD",X"44",X"4B",X"BC",X"00",X"0B",X"00",X"04",X"33",X"44",X"D7",X"BB",X"4B",X"CD",X"00",
		X"0B",X"00",X"0D",X"C7",X"BB",X"BC",X"BC",X"DC",X"D0",X"00",X"0B",X"00",X"D4",X"44",X"BB",X"B8",
		X"DD",X"8D",X"00",X"00",X"0B",X"D0",X"DC",X"BC",X"4C",X"DD",X"DD",X"D0",X"00",X"00",X"0C",X"BB",
		X"B7",X"BC",X"4D",X"DD",X"8D",X"D0",X"00",X"00",X"00",X"CC",X"BB",X"CC",X"48",X"DD",X"8D",X"CC",
		X"00",X"00",X"00",X"0D",X"DD",X"D4",X"C8",X"DD",X"C8",X"DD",X"00",X"00",X"00",X"00",X"84",X"CC",
		X"BD",X"DB",X"D8",X"DD",X"00",X"00",X"00",X"00",X"00",X"BB",X"BC",X"8D",X"D8",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"BB",X"BB",X"8D",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"DC",X"BB",X"8D",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DC",X"D0",X"00",X"00",X"00",X"00",X"97",X"57",
		X"90",X"00",X"A9",X"11",X"1A",X"00",X"09",X"91",X"60",X"00",X"00",X"A0",X"00",X"00",X"00",X"E5",
		X"09",X"00",X"90",X"00",X"00",X"A0",X"98",X"9F",X"97",X"00",X"70",X"00",X"0E",X"5A",X"81",X"88",
		X"15",X"00",X"00",X"0A",X"09",X"A8",X"88",X"89",X"57",X"00",X"00",X"07",X"E9",X"18",X"65",X"A0",
		X"00",X"00",X"90",X"00",X"5A",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"70",X"00",X"00",X"0E",
		X"0A",X"0E",X"00",X"A0",X"00",X"00",X"F0",X"00",X"A0",X"09",X"0F",X"0A",X"00",X"0A",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"90",X"0E",X"00",X"00",X"00",X"00",
		X"05",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"A0",X"00",X"0F",X"09",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"04",X"26",X"30",X"00",
		X"B0",X"00",X"00",X"00",X"00",X"00",X"36",X"42",X"30",X"00",X"B0",X"00",X"00",X"00",X"00",X"42",
		X"22",X"30",X"00",X"0C",X"BD",X"00",X"00",X"00",X"03",X"22",X"34",X"00",X"00",X"0C",X"BB",X"44",
		X"4D",X"C8",X"22",X"33",X"40",X"00",X"00",X"0D",X"CB",X"4B",X"B7",X"D4",X"43",X"34",X"00",X"0B",
		X"00",X"00",X"DC",X"DC",X"BC",X"BB",X"B7",X"CD",X"00",X"0B",X"00",X"00",X"0D",X"8D",X"D8",X"BB",
		X"B4",X"44",X"D0",X"0B",X"00",X"00",X"00",X"DD",X"DD",X"DC",X"4C",X"BC",X"D0",X"DB",X"00",X"00",
		X"00",X"DD",X"8D",X"DD",X"4C",X"B7",X"BB",X"BC",X"00",X"00",X"0C",X"CD",X"8D",X"D8",X"4C",X"CB",
		X"BC",X"C0",X"00",X"00",X"0D",X"D8",X"CD",X"D8",X"C4",X"DD",X"DD",X"00",X"00",X"00",X"0D",X"D8",
		X"DB",X"DD",X"BC",X"C4",X"80",X"00",X"00",X"00",X"00",X"D8",X"DD",X"8C",X"BB",X"B0",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"DD",X"8B",X"BB",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"8B",
		X"BC",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DC",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"97",X"57",X"90",X"0A",X"11",X"19",X"A0",X"00",X"61",X"99",X"00",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"90",X"09",X"05",X"E0",X"00",X"00",X"70",X"07",X"9F",X"98",X"90",X"A0",X"00",X"05",X"18",
		X"81",X"8A",X"5E",X"00",X"07",X"59",X"88",X"88",X"A9",X"0A",X"00",X"00",X"A5",X"68",X"19",X"E7",
		X"00",X"00",X"00",X"00",X"0A",X"50",X"00",X"90",X"00",X"00",X"00",X"70",X"07",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"0E",X"0A",X"0E",X"00",X"0A",X"0F",X"09",X"00",X"A0",X"00",X"F0",X"00",X"50",
		X"00",X"00",X"00",X"0A",X"00",X"90",X"00",X"00",X"00",X"0A",X"00",X"00",X"05",X"00",X"00",X"00",
		X"00",X"0E",X"00",X"A0",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"60",X"00",X"09",X"0F",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"09",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"05",X"05",X"00",X"05",X"95",X"00",X"00",X"90",X"00",X"09",
		X"79",X"00",X"0E",X"EE",X"00",X"05",X"55",X"00",X"00",X"70",X"00",X"00",X"05",X"05",X"00",X"00",
		X"00",X"05",X"95",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"19",X"79",X"10",X"00",X"01",
		X"A1",X"11",X"A1",X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"50",X"00",X"90",X"0A",X"00",X"00",
		X"00",X"00",X"A0",X"70",X"A0",X"00",X"00",X"00",X"7F",X"A9",X"89",X"AF",X"70",X"00",X"90",X"07",
		X"98",X"88",X"97",X"00",X"50",X"00",X"95",X"88",X"88",X"85",X"90",X"00",X"0A",X"05",X"8A",X"8A",
		X"85",X"0A",X"00",X"00",X"10",X"97",X"07",X"90",X"10",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0F",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"0F",X"0F",X"00",X"90",X"00",X"90",X"0E",X"00",X"00",X"A0",X"00",X"E0",X"0E",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"F0",X"F0",X"0E",X"00",X"00",X"00",X"F0",X"0E",X"00",X"90",X"E0",X"FE",X"00",X"00",X"A0",X"90",
		X"00",X"05",X"00",X"E0",X"E9",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"08",X"88",X"88",X"88",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"00",X"07",X"00",X"10",X"07",X"00",X"00",X"09",X"00",X"16",X"16",
		X"10",X"09",X"00",X"00",X"07",X"61",X"81",X"67",X"00",X"00",X"97",X"11",X"18",X"88",X"11",X"17",
		X"90",X"00",X"07",X"61",X"81",X"67",X"00",X"00",X"09",X"00",X"16",X"16",X"10",X"09",X"00",X"00",
		X"07",X"00",X"10",X"07",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"70",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"10",X"10",X"10",X"05",X"00",X"00",X"00",
		X"00",X"09",X"00",X"70",X"69",X"99",X"60",X"70",X"09",X"00",X"00",X"00",X"00",X"00",X"91",X"09",
		X"89",X"01",X"90",X"00",X"00",X"00",X"00",X"09",X"17",X"99",X"98",X"88",X"99",X"97",X"19",X"00",
		X"00",X"00",X"00",X"00",X"99",X"88",X"88",X"89",X"90",X"00",X"00",X"00",X"09",X"71",X"11",X"98",
		X"88",X"88",X"88",X"91",X"11",X"79",X"00",X"00",X"00",X"00",X"99",X"88",X"88",X"89",X"90",X"00",
		X"00",X"00",X"00",X"09",X"17",X"99",X"98",X"88",X"99",X"97",X"19",X"00",X"00",X"00",X"00",X"00",
		X"01",X"09",X"89",X"01",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"70",X"69",X"99",X"60",X"70",
		X"09",X"00",X"00",X"00",X"00",X"05",X"00",X"10",X"10",X"10",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"70",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"90",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"70",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"50",X"00",X"70",
		X"00",X"50",X"00",X"90",X"00",X"00",X"00",X"90",X"05",X"90",X"07",X"00",X"10",X"07",X"00",X"95",
		X"00",X"90",X"00",X"00",X"00",X"00",X"99",X"09",X"90",X"90",X"99",X"09",X"90",X"00",X"00",X"00",
		X"00",X"00",X"09",X"99",X"98",X"99",X"99",X"98",X"99",X"99",X"00",X"00",X"00",X"00",X"05",X"00",
		X"99",X"89",X"89",X"89",X"89",X"89",X"90",X"05",X"00",X"00",X"90",X"00",X"79",X"99",X"88",X"98",
		X"88",X"98",X"89",X"99",X"70",X"00",X"90",X"00",X"90",X"99",X"88",X"98",X"88",X"88",X"88",X"98",
		X"89",X"90",X"90",X"00",X"00",X"00",X"09",X"98",X"88",X"88",X"88",X"88",X"88",X"99",X"00",X"00",
		X"00",X"95",X"77",X"19",X"88",X"98",X"88",X"88",X"88",X"98",X"89",X"17",X"75",X"90",X"00",X"00",
		X"09",X"98",X"88",X"88",X"88",X"88",X"88",X"99",X"00",X"00",X"00",X"09",X"00",X"99",X"88",X"98",
		X"88",X"88",X"88",X"98",X"89",X"90",X"09",X"00",X"00",X"05",X"79",X"99",X"88",X"98",X"88",X"98",
		X"89",X"99",X"75",X"00",X"00",X"00",X"90",X"00",X"99",X"89",X"89",X"89",X"89",X"89",X"90",X"00",
		X"90",X"00",X"00",X"00",X"09",X"99",X"98",X"99",X"99",X"98",X"99",X"99",X"00",X"00",X"00",X"09",
		X"00",X"05",X"90",X"09",X"90",X"90",X"99",X"00",X"95",X"00",X"09",X"00",X"00",X"00",X"90",X"00",
		X"07",X"00",X"10",X"07",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"70",
		X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"A0",X"70",X"A0",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"0F",X"00",X"A0",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"0A",X"00",X"90",X"0A",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"0E",X"00",X"09",X"00",X"A0",X"0A",X"00",X"00",X"A0",X"00",X"0A",X"00",X"A0",X"09",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"A0",X"F0",X"00",X"90",X"00",X"F0",X"00",X"90",X"00",X"F0",
		X"A0",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"F0",X"00",X"F0",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"90",X"F0",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"F0",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0F",X"00",X"A9",X"5A",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"59",X"A0",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"09",X"00",X"00",X"00",
		X"00",X"F0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"F0",X"00",X"00",X"90",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"90",
		X"00",X"00",X"00",X"09",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"F0",X"00",X"A0",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"09",X"00",X"00",X"0A",X"00",X"00",X"00",X"0F",X"00",X"90",X"00",X"F0",X"00",X"90",
		X"0F",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"09",X"0A",X"00",X"0A",X"00",X"00",X"A0",X"00",
		X"0A",X"00",X"0A",X"09",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"0A",X"00",X"90",
		X"0A",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"0F",X"00",X"00",
		X"A0",X"0F",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"EE",
		X"EF",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"EE",X"EE",X"EF",X"FF",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"EE",X"EE",X"EF",X"FF",X"F0",X"00",X"E0",X"00",X"00",X"00",X"00",X"0E",X"EE",X"EE",
		X"EF",X"FF",X"F0",X"0E",X"F0",X"00",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"EF",X"FF",X"F8",X"E4",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"FF",X"FF",X"FF",X"40",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"EE",X"EF",X"FF",X"FF",X"F4",X"00",X"00",X"00",X"4E",X"EE",X"40",X"0F",X"EE",X"EE",
		X"FF",X"FF",X"40",X"00",X"00",X"00",X"09",X"88",X"E0",X"00",X"EE",X"EF",X"FF",X"F4",X"00",X"00",
		X"00",X"00",X"EE",X"EE",X"E0",X"00",X"F8",X"8F",X"F4",X"00",X"00",X"00",X"00",X"04",X"EF",X"FF",
		X"E0",X"00",X"EE",X"8F",X"40",X"00",X"00",X"00",X"00",X"4E",X"00",X"0F",X"FE",X"EE",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"EE",X"F0",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"0F",X"EE",X"F0",X"00",X"00",X"09",X"A0",X"00",X"00",X"00",X"0F",X"EE",X"F0",X"00",
		X"FA",X"9A",X"FF",X"00",X"00",X"00",X"0F",X"EE",X"F0",X"0F",X"88",X"88",X"8E",X"E0",X"00",X"00",
		X"0F",X"EF",X"F0",X"04",X"58",X"87",X"8A",X"EF",X"00",X"00",X"0F",X"EF",X"40",X"4F",X"8E",X"F8",
		X"89",X"CF",X"40",X"00",X"FE",X"FF",X"00",X"A9",X"9F",X"82",X"56",X"F3",X"F4",X"3F",X"2F",X"F0",
		X"00",X"95",X"F4",X"99",X"E3",X"FF",X"33",X"33",X"FF",X"00",X"00",X"5A",X"A9",X"AF",X"00",X"0F",
		X"FF",X"FF",X"40",X"00",X"00",X"5A",X"AF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"EE",X"F0",X"00",X"00",X"00",X"00",X"0F",X"EE",
		X"F0",X"00",X"00",X"00",X"00",X"0F",X"EE",X"F0",X"00",X"00",X"00",X"00",X"0F",X"EE",X"F0",X"00",
		X"00",X"00",X"00",X"0F",X"EF",X"F0",X"00",X"00",X"00",X"00",X"0F",X"EF",X"F0",X"00",X"00",X"00",
		X"00",X"0F",X"EF",X"40",X"00",X"00",X"00",X"00",X"0E",X"FF",X"00",X"00",X"00",X"90",X"00",X"FE",
		X"F4",X"00",X"00",X"A9",X"A0",X"0F",X"EF",X"F0",X"00",X"09",X"AF",X"9F",X"EE",X"FF",X"00",X"00",
		X"88",X"88",X"8E",X"AE",X"20",X"00",X"00",X"58",X"87",X"83",X"9B",X"F0",X"00",X"00",X"A8",X"38",
		X"32",X"6F",X"00",X"00",X"00",X"5E",X"83",X"99",X"F0",X"00",X"00",X"00",X"5E",X"49",X"AF",X"00",
		X"00",X"00",X"00",X"95",X"AA",X"F0",X"00",X"00",X"00",X"00",X"09",X"9A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A9",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"80",X"00",X"00",
		X"00",X"08",X"88",X"88",X"88",X"00",X"00",X"08",X"88",X"08",X"88",X"88",X"80",X"00",X"88",X"80",
		X"08",X"88",X"88",X"80",X"00",X"08",X"88",X"88",X"00",X"88",X"80",X"00",X"88",X"80",X"88",X"08",
		X"88",X"00",X"08",X"00",X"88",X"88",X"88",X"80",X"00",X"00",X"88",X"08",X"08",X"80",X"00",X"00",
		X"00",X"08",X"80",X"00",X"00",X"00",X"00",X"FE",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FE",X"EF",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"FE",X"EF",X"00",X"00",X"00",
		X"00",X"A9",X"00",X"00",X"00",X"FE",X"EF",X"00",X"00",X"00",X"0F",X"FA",X"9A",X"F0",X"00",X"FF",
		X"EF",X"00",X"00",X"00",X"EE",X"88",X"88",X"8F",X"00",X"4F",X"EF",X"00",X"00",X"0F",X"EA",X"87",
		X"88",X"54",X"00",X"0F",X"FE",X"F0",X"00",X"4F",X"C9",X"88",X"FE",X"8F",X"40",X"00",X"FF",X"2F",
		X"34",X"F3",X"F6",X"52",X"8F",X"99",X"A0",X"00",X"0F",X"F3",X"33",X"3F",X"F3",X"E9",X"94",X"F5",
		X"90",X"00",X"00",X"4F",X"FF",X"FF",X"00",X"0F",X"A9",X"AA",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"AA",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"FE",X"EF",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"EF",X"00",X"00",X"00",X"00",X"00",X"FE",X"EF",X"00",X"00",X"00",X"00",X"00",X"FE",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"EF",X"00",X"00",X"00",X"00",X"00",X"FF",X"EF",X"00",X"00",
		X"00",X"00",X"00",X"4F",X"EF",X"00",X"00",X"00",X"00",X"00",X"0F",X"FE",X"00",X"00",X"00",X"00",
		X"00",X"04",X"FE",X"F0",X"00",X"90",X"00",X"00",X"00",X"FF",X"EF",X"00",X"A9",X"A0",X"00",X"00",
		X"0F",X"FE",X"EF",X"9F",X"A9",X"00",X"00",X"00",X"2E",X"AE",X"88",X"88",X"80",X"00",X"00",X"FB",
		X"93",X"87",X"88",X"50",X"00",X"00",X"0F",X"62",X"38",X"38",X"A0",X"00",X"00",X"00",X"F9",X"93",
		X"8E",X"50",X"00",X"00",X"00",X"0F",X"A9",X"4E",X"50",X"00",X"00",X"00",X"00",X"FA",X"A5",X"90",
		X"00",X"00",X"00",X"00",X"0A",X"99",X"00",X"00",X"00",X"00",X"00",X"A9",X"A0",X"00",X"00",X"88",
		X"88",X"80",X"00",X"00",X"00",X"08",X"88",X"88",X"88",X"00",X"00",X"00",X"88",X"88",X"88",X"08",
		X"88",X"00",X"00",X"88",X"88",X"88",X"00",X"88",X"80",X"00",X"88",X"80",X"08",X"88",X"88",X"00",
		X"00",X"08",X"88",X"08",X"80",X"88",X"80",X"00",X"00",X"88",X"88",X"88",X"80",X"08",X"00",X"00",
		X"00",X"88",X"08",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"0F",
		X"EE",X"F0",X"00",X"00",X"0F",X"EE",X"F0",X"00",X"00",X"0F",X"EE",X"F0",X"00",X"00",X"0F",X"EE",
		X"F0",X"00",X"00",X"0F",X"E3",X"F0",X"00",X"00",X"04",X"EF",X"F0",X"00",X"00",X"00",X"EF",X"F0",
		X"00",X"00",X"00",X"EF",X"F0",X"00",X"00",X"00",X"EF",X"F0",X"00",X"00",X"00",X"EF",X"F0",X"AF",
		X"00",X"4F",X"EF",X"F0",X"09",X"AF",X"FF",X"2E",X"F0",X"00",X"9E",X"FE",X"9B",X"F0",X"00",X"A8",
		X"88",X"95",X"F0",X"00",X"0F",X"78",X"F6",X"F0",X"00",X"0F",X"FF",X"9E",X"30",X"00",X"00",X"5F",
		X"A9",X"00",X"00",X"00",X"A5",X"EA",X"00",X"00",X"00",X"0A",X"99",X"F0",X"FE",X"EF",X"00",X"00",
		X"00",X"FE",X"EF",X"00",X"00",X"00",X"FE",X"EF",X"00",X"00",X"00",X"FE",X"EF",X"00",X"00",X"00",
		X"F3",X"EF",X"00",X"00",X"00",X"FF",X"E4",X"00",X"00",X"00",X"FF",X"E0",X"00",X"00",X"00",X"FF",
		X"E0",X"00",X"00",X"00",X"FF",X"E0",X"00",X"00",X"00",X"FF",X"E0",X"00",X"00",X"00",X"FF",X"EF",
		X"40",X"0F",X"A0",X"FE",X"2F",X"FF",X"A9",X"00",X"FB",X"9E",X"FE",X"90",X"00",X"F5",X"98",X"88",
		X"A0",X"00",X"F6",X"F8",X"7F",X"00",X"00",X"3E",X"9F",X"FF",X"00",X"00",X"09",X"AF",X"50",X"00",
		X"00",X"0A",X"E5",X"A0",X"00",X"00",X"F9",X"9A",X"00",X"00",X"00",X"0A",X"A9",X"AA",X"00",X"00",
		X"00",X"A9",X"55",X"99",X"A0",X"00",X"00",X"0A",X"55",X"99",X"9A",X"00",X"00",X"00",X"A9",X"55",
		X"59",X"A0",X"00",X"00",X"0A",X"A9",X"99",X"9A",X"00",X"00",X"0A",X"9A",X"00",X"00",X"00",X"A9",
		X"59",X"90",X"00",X"0A",X"A9",X"95",X"9A",X"00",X"0A",X"A9",X"95",X"99",X"00",X"0A",X"AA",X"99",
		X"9A",X"00",X"00",X"AA",X"AA",X"90",X"00",X"00",X"0A",X"AA",X"00",X"00",X"00",X"0A",X"8A",X"00",
		X"00",X"00",X"A8",X"98",X"90",X"00",X"0A",X"8A",X"98",X"99",X"00",X"0A",X"8A",X"98",X"99",X"00",
		X"0A",X"AA",X"98",X"9A",X"00",X"00",X"AA",X"9A",X"90",X"00",X"00",X"0A",X"AA",X"00",X"00",X"00",
		X"0F",X"EF",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A8",X"A9",
		X"00",X"00",X"09",X"88",X"88",X"89",X"00",X"0A",X"8A",X"98",X"99",X"00",X"0A",X"8A",X"98",X"99",
		X"00",X"0A",X"8A",X"98",X"99",X"00",X"0A",X"8A",X"98",X"99",X"00",X"0A",X"AA",X"98",X"9A",X"00",
		X"00",X"AA",X"9A",X"90",X"00",X"00",X"0A",X"AA",X"00",X"00",X"00",X"0F",X"EF",X"00",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"A9",X"00",
		X"00",X"09",X"88",X"88",X"89",X"00",X"0A",X"89",X"98",X"99",X"00",X"0A",X"8A",X"98",X"99",X"00",
		X"0A",X"8A",X"98",X"99",X"00",X"0A",X"8A",X"98",X"99",X"00",X"0A",X"8A",X"98",X"99",X"00",X"0A",
		X"8A",X"98",X"99",X"00",X"0A",X"8A",X"98",X"99",X"00",X"0A",X"AA",X"98",X"9A",X"00",X"00",X"AA",
		X"9A",X"90",X"00",X"00",X"0A",X"AA",X"00",X"00",X"00",X"FF",X"EF",X"00",X"00",X"00",X"FE",X"EF",
		X"00",X"00",X"00",X"0F",X"E0",X"00",X"00",X"00",X"0F",X"EF",X"00",X"00",X"00",X"0F",X"E0",X"00",
		X"00",X"00",X"FF",X"E0",X"00",X"00",X"00",X"0F",X"E0",X"00",X"00",X"00",X"0F",X"90",X"00",X"00",
		X"00",X"0F",X"E0",X"00",X"00",X"00",X"0F",X"9F",X"00",X"00",X"00",X"0E",X"90",X"00",X"00",X"00",
		X"0E",X"90",X"00",X"00",X"00",X"0F",X"90",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"9A",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"90",
		X"00",X"09",X"99",X"00",X"00",X"00",X"09",X"99",X"00",X"0A",X"9A",X"00",X"00",X"00",X"00",X"A9",
		X"A0",X"0A",X"9A",X"00",X"A9",X"00",X"00",X"09",X"9A",X"09",X"9A",X"00",X"99",X"A0",X"99",X"0A",
		X"88",X"88",X"8A",X"09",X"9A",X"00",X"09",X"98",X"8E",X"6E",X"88",X"A9",X"A0",X"00",X"00",X"A9",
		X"A8",X"E1",X"88",X"9A",X"00",X"00",X"00",X"0A",X"A9",X"A8",X"89",X"90",X"00",X"00",X"00",X"00",
		X"AA",X"98",X"99",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"E4",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"E0",X"90",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"EE",X"90",X"00",X"00",X"00",X"00",X"00",X"FE",X"99",X"90",X"00",X"00",X"00",X"00",X"00",
		X"FB",X"9A",X"A0",X"00",X"00",X"00",X"00",X"00",X"F5",X"98",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"F6",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"FE",X"9F",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"09",X"A5",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"5A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F9",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"A9",X"AA",X"00",X"00",X"00",X"A9",X"95",
		X"59",X"A0",X"00",X"0A",X"99",X"95",X"5A",X"00",X"00",X"A9",X"55",X"59",X"A0",X"00",X"0A",X"99",
		X"99",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"89",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8A",X"9A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"89",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"88",X"80",X"00",X"00",X"00",X"00",X"09",X"AA",X"AA",X"9A",X"8E",
		X"19",X"8A",X"9A",X"AA",X"99",X"00",X"99",X"99",X"99",X"88",X"86",X"E7",X"88",X"89",X"99",X"99",
		X"90",X"89",X"9A",X"AA",X"A9",X"88",X"88",X"89",X"AA",X"AA",X"99",X"00",X"08",X"88",X"88",X"88",
		X"89",X"89",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"8A",X"89",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"8A",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"89",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"9A",X"00",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"00",X"A9",X"9A",X"00",X"00",X"00",X"0A",X"99",X"9A",X"00",X"00",X"09",X"9A",
		X"A8",X"00",X"00",X"00",X"08",X"A9",X"99",X"A9",X"88",X"88",X"89",X"80",X"00",X"00",X"00",X"00",
		X"88",X"AA",X"98",X"8E",X"6E",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"9A",X"87",X"91",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"9A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"89",X"A8",X"99",X"99",X"9A",X"A0",X"00",X"00",X"00",X"00",X"99",X"9A",
		X"80",X"88",X"AA",X"99",X"9A",X"00",X"00",X"00",X"09",X"99",X"A8",X"00",X"00",X"88",X"8A",X"A0",
		X"00",X"00",X"00",X"0A",X"9A",X"80",X"00",X"00",X"00",X"08",X"80",X"00",X"00",X"00",X"08",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"99",X"A0",X"00",X"00",X"00",X"0A",X"A0",X"00",X"00",X"00",X"08",
		X"AA",X"89",X"00",X"00",X"0A",X"A9",X"9A",X"00",X"00",X"00",X"00",X"8A",X"88",X"88",X"AA",X"A9",
		X"99",X"A8",X"00",X"00",X"00",X"00",X"08",X"89",X"7E",X"88",X"9A",X"A8",X"80",X"00",X"00",X"00",
		X"00",X"09",X"81",X"E6",X"8A",X"98",X"80",X"00",X"00",X"00",X"00",X"0A",X"98",X"88",X"88",X"88",
		X"80",X"00",X"00",X"00",X"00",X"0A",X"99",X"99",X"98",X"A9",X"89",X"00",X"00",X"00",X"00",X"0A",
		X"99",X"9A",X"A8",X"80",X"8A",X"AA",X"90",X"00",X"00",X"00",X"08",X"9A",X"A8",X"80",X"00",X"08",
		X"A9",X"99",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"8A",X"9A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"80",X"00",X"00",X"00",X"E4",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"E0",X"EE",X"40",X"00",X"0F",X"EE",X"EF",X"40",X"00",
		X"00",X"00",X"F9",X"8E",X"F0",X"00",X"EE",X"EE",X"EF",X"FF",X"00",X"00",X"00",X"FF",X"EE",X"F0",
		X"0F",X"EE",X"EE",X"EF",X"FF",X"40",X"00",X"00",X"0E",X"EE",X"00",X"0E",X"EE",X"EE",X"EF",X"FF",
		X"F0",X"00",X"00",X"0F",X"F0",X"00",X"0E",X"EE",X"EE",X"EF",X"FF",X"F0",X"00",X"00",X"0E",X"FF",
		X"00",X"0E",X"EE",X"EE",X"EF",X"FF",X"F0",X"00",X"00",X"00",X"EF",X"F0",X"8E",X"EE",X"EE",X"FF",
		X"FF",X"F0",X"00",X"00",X"00",X"0E",X"FF",X"4E",X"EE",X"EF",X"FF",X"FF",X"F0",X"00",X"00",X"00",
		X"00",X"FF",X"4F",X"EE",X"FF",X"FF",X"FF",X"40",X"00",X"00",X"00",X"00",X"00",X"4F",X"FF",X"FF",
		X"FF",X"F4",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"FF",X"FF",X"FF",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"FF",X"FE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"4F",X"FE",X"EF",X"F0",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"05",
		X"59",X"AF",X"40",X"98",X"00",X"00",X"00",X"00",X"79",X"E3",X"88",X"A9",X"A4",X"00",X"00",X"00",
		X"05",X"2A",X"88",X"58",X"A9",X"AE",X"00",X"00",X"00",X"09",X"9A",X"9F",X"8A",X"9E",X"FE",X"00",
		X"00",X"00",X"09",X"4A",X"A9",X"E9",X"EE",X"FE",X"00",X"00",X"00",X"0A",X"00",X"FE",X"59",X"EF",
		X"F3",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"3F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"43",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"EF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"F4",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EF",X"F3",X"0F",X"EF",X"F0",X"00",X"00",X"00",X"00",X"4E",X"FF",
		X"FE",X"FF",X"F0",X"00",X"00",X"00",X"00",X"04",X"FF",X"FF",X"FF",X"40",X"00",X"00",X"00",X"00",
		X"00",X"44",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"A9",X"00",X"0F",X"EE",X"F0",X"00",X"05",X"5A",X"84",X"A9",X"A4",X"0F",X"EE",X"F0",
		X"00",X"79",X"E8",X"58",X"AA",X"AE",X"0F",X"EE",X"F0",X"05",X"2A",X"88",X"88",X"9E",X"FE",X"0F",
		X"EE",X"F0",X"09",X"9A",X"9F",X"AA",X"9E",X"F3",X"0F",X"EF",X"F0",X"09",X"4A",X"A9",X"79",X"EE",
		X"F0",X"0F",X"EF",X"40",X"0A",X"00",X"40",X"49",X"EF",X"30",X"0E",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"4E",X"FF",X"EF",X"F0",X"00",X"00",X"00",X"00",X"00",X"04",X"3F",X"FF",X"00",X"00",X"20",
		X"49",X"4E",X"46",X"45",X"52",X"4E",X"4F",X"20",X"2D",X"20",X"43",X"4F",X"50",X"59",X"52",X"49",
		X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",X"38",X"34",X"20",X"57",X"49",X"4C",
		X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",
		X"53",X"20",X"49",X"4E",X"43",X"2E",X"00",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"88",X"08",
		X"08",X"80",X"00",X"00",X"08",X"80",X"88",X"88",X"88",X"80",X"00",X"00",X"08",X"88",X"08",X"80",
		X"88",X"00",X"00",X"08",X"88",X"88",X"00",X"88",X"80",X"00",X"88",X"88",X"08",X"88",X"88",X"80",
		X"00",X"08",X"80",X"08",X"88",X"88",X"80",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",
		X"00",X"88",X"88",X"80",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"90",X"4F",X"A9",X"55",X"00",X"00",X"00",X"00",X"04",X"A9",X"A8",X"83",X"E9",X"70",X"00",
		X"00",X"00",X"0E",X"A9",X"A8",X"58",X"8A",X"25",X"00",X"00",X"00",X"0E",X"FE",X"9A",X"8F",X"9A",
		X"99",X"00",X"00",X"00",X"0E",X"FE",X"E9",X"E9",X"AA",X"49",X"00",X"00",X"00",X"03",X"FF",X"E9",
		X"5E",X"F0",X"0A",X"00",X"00",X"00",X"00",X"FF",X"3C",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"FF",X"E0",X"00",X"00",X"00",
		X"00",X"FF",X"EF",X"03",X"FF",X"E0",X"00",X"00",X"00",X"00",X"FF",X"FE",X"FF",X"FE",X"40",X"00",
		X"00",X"00",X"00",X"4F",X"FF",X"FF",X"F4",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"F4",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"FE",X"EF",
		X"00",X"09",X"A4",X"00",X"00",X"00",X"00",X"FE",X"EF",X"04",X"A9",X"A4",X"8A",X"55",X"00",X"00",
		X"FE",X"EF",X"0E",X"AA",X"A8",X"58",X"E9",X"70",X"00",X"FE",X"EF",X"0E",X"FE",X"98",X"88",X"8A",
		X"25",X"00",X"FF",X"EF",X"03",X"FE",X"9A",X"AF",X"9A",X"99",X"00",X"4F",X"EF",X"00",X"FE",X"E9",
		X"79",X"AA",X"49",X"00",X"0F",X"FE",X"00",X"3F",X"E9",X"40",X"40",X"0A",X"00",X"00",X"FF",X"EF",
		X"FE",X"40",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"34",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"88",X"08",X"08",X"80",X"00",X"00",X"88",X"88",
		X"88",X"80",X"88",X"00",X"08",X"80",X"88",X"08",X"88",X"00",X"00",X"88",X"80",X"08",X"88",X"88",
		X"00",X"00",X"88",X"88",X"88",X"08",X"88",X"80",X"00",X"88",X"88",X"88",X"00",X"88",X"00",X"00",
		X"08",X"88",X"88",X"88",X"80",X"00",X"00",X"00",X"88",X"88",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"07",X"00",X"09",X"79",
		X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"05",X"75",X"09",X"70",X"00",X"90",X"00",
		X"00",X"07",X"00",X"91",X"55",X"15",X"51",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"75",
		X"75",X"75",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"55",X"57",X"77",X"55",X"59",X"00",X"00",
		X"00",X"01",X"77",X"17",X"71",X"77",X"17",X"71",X"77",X"17",X"71",X"00",X"00",X"00",X"09",X"55",
		X"57",X"77",X"55",X"59",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"75",X"75",X"75",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"91",X"55",X"15",X"51",X"90",X"07",X"00",X"00",X"00",X"90",X"00",
		X"79",X"05",X"75",X"09",X"70",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"09",X"79",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"07",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"10",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"09",X"79",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"19",X"05",X"15",X"09",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"97",
		X"55",X"75",X"57",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"75",X"75",X"75",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"55",X"51",X"11",X"55",X"59",X"00",X"00",X"00",X"70",X"71",X"77",
		X"17",X"71",X"71",X"77",X"17",X"71",X"70",X"70",X"00",X"00",X"09",X"55",X"51",X"11",X"55",X"59",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"75",X"75",X"75",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"97",X"55",X"75",X"57",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"05",X"15",X"09",
		X"10",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"09",X"79",X"00",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"10",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"09",X"19",X"00",X"01",X"00",X"00",X"00",X"00",X"79",X"05",X"75",X"09",
		X"70",X"00",X"00",X"00",X"00",X"97",X"55",X"75",X"57",X"90",X"00",X"00",X"00",X"00",X"05",X"15",
		X"15",X"15",X"00",X"00",X"00",X"00",X"09",X"55",X"57",X"77",X"55",X"59",X"00",X"00",X"17",X"71",
		X"77",X"17",X"77",X"17",X"71",X"77",X"10",X"00",X"09",X"55",X"57",X"77",X"55",X"59",X"00",X"00",
		X"00",X"00",X"05",X"15",X"15",X"15",X"00",X"00",X"00",X"00",X"00",X"97",X"55",X"75",X"57",X"90",
		X"00",X"00",X"00",X"00",X"79",X"05",X"75",X"09",X"70",X"00",X"00",X"00",X"01",X"00",X"09",X"19",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"06",X"00",X"03",
		X"63",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"63",X"02",X"62",X"03",X"60",X"00",X"20",
		X"00",X"00",X"06",X"00",X"31",X"22",X"12",X"21",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"62",X"62",X"62",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"22",X"26",X"66",X"22",X"23",X"00",
		X"00",X"00",X"01",X"66",X"16",X"61",X"66",X"16",X"61",X"66",X"16",X"61",X"00",X"00",X"00",X"03",
		X"22",X"26",X"66",X"22",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"62",X"62",X"62",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"22",X"12",X"21",X"30",X"06",X"00",X"00",X"00",X"20",
		X"00",X"63",X"02",X"62",X"03",X"60",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"03",X"63",X"00",
		X"06",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"06",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"10",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"03",X"63",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"13",X"02",X"12",X"03",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"36",X"22",X"62",X"26",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"62",X"62",X"62",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"22",X"21",X"11",X"22",X"23",X"00",X"00",X"00",X"60",X"61",
		X"66",X"16",X"61",X"61",X"66",X"16",X"61",X"60",X"60",X"00",X"00",X"03",X"22",X"21",X"11",X"22",
		X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"62",X"62",X"62",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"36",X"22",X"62",X"26",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"02",X"12",
		X"03",X"10",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"03",X"63",X"00",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"10",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"03",X"13",X"00",X"01",X"00",X"00",X"00",X"00",X"63",X"02",X"62",
		X"03",X"60",X"00",X"00",X"00",X"00",X"36",X"22",X"62",X"26",X"30",X"00",X"00",X"00",X"00",X"02",
		X"12",X"12",X"12",X"00",X"00",X"00",X"00",X"03",X"22",X"26",X"66",X"22",X"23",X"00",X"00",X"16",
		X"61",X"66",X"16",X"66",X"16",X"61",X"66",X"10",X"00",X"03",X"22",X"26",X"66",X"22",X"23",X"00",
		X"00",X"00",X"00",X"02",X"12",X"12",X"12",X"00",X"00",X"00",X"00",X"00",X"36",X"22",X"62",X"26",
		X"30",X"00",X"00",X"00",X"00",X"63",X"02",X"62",X"03",X"60",X"00",X"00",X"00",X"01",X"00",X"03",
		X"13",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"11",X"17",X"77",X"55",X"59",X"99",X"10",X"11",X"17",X"77",X"55",X"59",X"99",X"10",X"11",X"17",
		X"77",X"55",X"59",X"99",X"10",X"11",X"17",X"77",X"55",X"59",X"99",X"10",X"11",X"17",X"77",X"55",
		X"59",X"99",X"10",X"11",X"17",X"77",X"55",X"59",X"99",X"10",X"11",X"17",X"77",X"55",X"59",X"99",
		X"10",X"11",X"17",X"77",X"55",X"59",X"99",X"10",X"11",X"17",X"77",X"55",X"59",X"99",X"10",X"11",
		X"17",X"77",X"55",X"59",X"99",X"10",X"11",X"17",X"77",X"55",X"59",X"99",X"10",X"11",X"17",X"77",
		X"55",X"59",X"99",X"10",X"11",X"17",X"77",X"55",X"59",X"99",X"10",X"11",X"17",X"77",X"55",X"59",
		X"99",X"10",X"11",X"17",X"77",X"55",X"59",X"99",X"10",X"11",X"17",X"77",X"55",X"59",X"99",X"10",
		X"11",X"17",X"77",X"55",X"59",X"99",X"10",X"11",X"17",X"77",X"55",X"59",X"99",X"10",X"11",X"17",
		X"77",X"55",X"59",X"99",X"10",X"11",X"17",X"77",X"55",X"59",X"99",X"10",X"11",X"17",X"77",X"55",
		X"59",X"99",X"10",X"01",X"17",X"77",X"55",X"59",X"99",X"00",X"00",X"07",X"77",X"55",X"59",X"00",
		X"00",X"00",X"00",X"77",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"77",
		X"75",X"55",X"99",X"91",X"11",X"70",X"77",X"75",X"55",X"99",X"91",X"11",X"70",X"77",X"75",X"55",
		X"99",X"91",X"11",X"70",X"77",X"75",X"55",X"99",X"91",X"11",X"70",X"77",X"75",X"55",X"99",X"91",
		X"11",X"70",X"77",X"75",X"55",X"99",X"91",X"11",X"70",X"77",X"75",X"55",X"99",X"91",X"11",X"70",
		X"77",X"75",X"55",X"99",X"91",X"11",X"70",X"77",X"75",X"55",X"99",X"91",X"11",X"70",X"77",X"75",
		X"55",X"99",X"91",X"11",X"70",X"77",X"75",X"55",X"99",X"91",X"11",X"70",X"77",X"75",X"55",X"99",
		X"91",X"11",X"70",X"77",X"75",X"55",X"99",X"91",X"11",X"70",X"77",X"75",X"55",X"99",X"91",X"11",
		X"70",X"77",X"75",X"55",X"99",X"91",X"11",X"70",X"77",X"75",X"55",X"99",X"91",X"11",X"70",X"77",
		X"75",X"55",X"99",X"91",X"11",X"70",X"77",X"75",X"55",X"99",X"91",X"11",X"70",X"77",X"75",X"55",
		X"99",X"91",X"11",X"70",X"77",X"75",X"55",X"99",X"91",X"11",X"70",X"77",X"75",X"55",X"99",X"91",
		X"11",X"70",X"07",X"75",X"55",X"99",X"91",X"11",X"00",X"00",X"05",X"55",X"99",X"91",X"00",X"00",
		X"00",X"00",X"55",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"55",X"59",
		X"99",X"11",X"17",X"77",X"50",X"55",X"59",X"99",X"11",X"17",X"77",X"50",X"55",X"59",X"99",X"11",
		X"17",X"77",X"50",X"55",X"59",X"99",X"11",X"17",X"77",X"50",X"55",X"59",X"99",X"11",X"17",X"77",
		X"50",X"55",X"59",X"99",X"11",X"17",X"77",X"50",X"55",X"59",X"99",X"11",X"17",X"77",X"50",X"55",
		X"59",X"99",X"11",X"17",X"77",X"50",X"55",X"59",X"99",X"11",X"17",X"77",X"50",X"55",X"59",X"99",
		X"11",X"17",X"77",X"50",X"55",X"59",X"99",X"11",X"17",X"77",X"50",X"55",X"59",X"99",X"11",X"17",
		X"77",X"50",X"55",X"59",X"99",X"11",X"17",X"77",X"50",X"55",X"59",X"99",X"11",X"17",X"77",X"50",
		X"55",X"59",X"99",X"11",X"17",X"77",X"50",X"55",X"59",X"99",X"11",X"17",X"77",X"50",X"55",X"59",
		X"99",X"11",X"17",X"77",X"50",X"55",X"59",X"99",X"11",X"17",X"77",X"50",X"55",X"59",X"99",X"11",
		X"17",X"77",X"50",X"55",X"59",X"99",X"11",X"17",X"77",X"50",X"55",X"59",X"99",X"11",X"17",X"77",
		X"50",X"05",X"59",X"99",X"11",X"17",X"77",X"00",X"00",X"09",X"99",X"11",X"17",X"00",X"00",X"00",
		X"00",X"99",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"99",X"91",X"11",
		X"77",X"75",X"55",X"90",X"99",X"91",X"11",X"77",X"75",X"55",X"90",X"99",X"91",X"11",X"77",X"75",
		X"55",X"90",X"99",X"91",X"11",X"77",X"75",X"55",X"90",X"99",X"91",X"11",X"77",X"75",X"55",X"90",
		X"99",X"91",X"11",X"77",X"75",X"55",X"90",X"99",X"91",X"11",X"77",X"75",X"55",X"90",X"99",X"91",
		X"11",X"77",X"75",X"55",X"90",X"99",X"91",X"11",X"77",X"75",X"55",X"90",X"99",X"91",X"11",X"77",
		X"75",X"55",X"90",X"99",X"91",X"11",X"77",X"75",X"55",X"90",X"99",X"91",X"11",X"77",X"75",X"55",
		X"90",X"99",X"91",X"11",X"77",X"75",X"55",X"90",X"99",X"91",X"11",X"77",X"75",X"55",X"90",X"99",
		X"91",X"11",X"77",X"75",X"55",X"90",X"99",X"91",X"11",X"77",X"75",X"55",X"90",X"99",X"91",X"11",
		X"77",X"75",X"55",X"90",X"99",X"91",X"11",X"77",X"75",X"55",X"90",X"99",X"91",X"11",X"77",X"75",
		X"55",X"90",X"99",X"91",X"11",X"77",X"75",X"55",X"90",X"99",X"91",X"11",X"77",X"75",X"55",X"90",
		X"09",X"91",X"11",X"77",X"75",X"55",X"00",X"00",X"01",X"11",X"77",X"75",X"00",X"00",X"00",X"00",
		X"11",X"77",X"70",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"80",X"00",X"00",X"00",X"08",X"88",X"88",X"88",X"00",
		X"00",X"08",X"88",X"88",X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"80",X"08",
		X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"08",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"88",
		X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"05",X"75",X"00",X"00",X"00",X"00",X"00",X"97",
		X"99",X"00",X"00",X"00",X"00",X"0A",X"99",X"59",X"00",X"00",X"00",X"00",X"A5",X"57",X"70",X"00",
		X"00",X"00",X"00",X"57",X"10",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"00",X"00",X"00",
		X"00",X"00",X"05",X"99",X"00",X"00",X"00",X"00",X"00",X"9A",X"59",X"00",X"00",X"00",X"00",X"09",
		X"57",X"79",X"00",X"00",X"00",X"00",X"A7",X"79",X"50",X"00",X"00",X"00",X"00",X"95",X"90",X"A0",
		X"00",X"00",X"00",X"00",X"0A",X"9A",X"00",X"00",X"00",X"00",X"95",X"79",X"00",X"00",X"00",X"0A",
		X"79",X"99",X"00",X"00",X"00",X"A9",X"55",X"50",X"00",X"00",X"00",X"95",X"70",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"00",X"00",X"05",X"75",X"00",X"00",X"00",
		X"09",X"97",X"90",X"00",X"00",X"09",X"59",X"9A",X"00",X"00",X"00",X"77",X"55",X"A0",X"00",X"00",
		X"00",X"17",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"09",X"70",X"00",X"00",X"00",X"09",X"95",X"00",X"00",X"00",X"09",X"5A",X"90",X"00",X"00",X"09",
		X"77",X"59",X"00",X"00",X"00",X"59",X"77",X"A0",X"00",X"00",X"00",X"95",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"0A",X"9A",X"00",X"00",X"09",X"75",X"90",X"00",
		X"09",X"99",X"7A",X"00",X"00",X"55",X"59",X"A0",X"00",X"00",X"75",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"57",X"10",X"00",X"00",X"00",X"A5",X"57",X"70",X"00",X"00",X"0A",X"99",X"59",
		X"00",X"00",X"00",X"97",X"99",X"00",X"00",X"00",X"05",X"75",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"90",X"00",
		X"00",X"00",X"A7",X"79",X"50",X"00",X"00",X"09",X"57",X"79",X"00",X"00",X"00",X"9A",X"59",X"00",
		X"00",X"00",X"05",X"99",X"00",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"70",X"00",X"00",X"A9",X"55",X"50",X"00",X"0A",X"79",
		X"99",X"00",X"00",X"95",X"79",X"00",X"00",X"0A",X"9A",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"17",X"50",X"00",X"00",X"00",X"00",X"77",X"55",X"A0",X"00",X"00",X"00",X"09",X"59",X"9A",
		X"00",X"00",X"00",X"00",X"09",X"97",X"90",X"00",X"00",X"00",X"00",X"05",X"75",X"00",X"00",X"00",
		X"00",X"00",X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"95",X"90",X"00",X"00",X"00",
		X"00",X"59",X"77",X"A0",X"00",X"00",X"00",X"09",X"77",X"59",X"00",X"00",X"00",X"00",X"09",X"5A",
		X"90",X"00",X"00",X"00",X"00",X"09",X"95",X"00",X"00",X"00",X"00",X"00",X"09",X"70",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"75",X"90",X"00",X"00",X"00",X"55",X"59",X"A0",X"00",X"00",X"09",
		X"99",X"7A",X"00",X"00",X"00",X"09",X"75",X"90",X"00",X"00",X"00",X"0A",X"9A",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"CC",X"BB",X"00",X"00",X"00",X"0B",X"CB",X"3B",X"B0",X"00",
		X"00",X"CC",X"BB",X"3B",X"B0",X"00",X"0C",X"BC",X"BC",X"CB",X"B0",X"00",X"BB",X"CC",X"CB",X"BB",
		X"00",X"0B",X"BC",X"0C",X"BB",X"CC",X"C0",X"0B",X"C0",X"0C",X"BB",X"CC",X"C0",X"00",X"B0",X"0C",
		X"BB",X"3B",X"B0",X"00",X"00",X"0B",X"CC",X"0B",X"B0",X"00",X"00",X"0B",X"B0",X"0B",X"C0",X"00",
		X"00",X"CB",X"B0",X"0B",X"B0",X"00",X"0C",X"BB",X"C0",X"0B",X"B0",X"00",X"0B",X"BC",X"00",X"CB",
		X"B0",X"00",X"00",X"00",X"0C",X"BB",X"C0",X"00",X"00",X"00",X"0B",X"BC",X"00",X"00",X"00",X"00",
		X"0C",X"BB",X"00",X"00",X"00",X"00",X"00",X"CB",X"3B",X"B0",X"00",X"00",X"0C",X"B3",X"CB",X"33",
		X"BB",X"00",X"BB",X"0B",X"CB",X"BB",X"C3",X"BB",X"00",X"BB",X"CB",X"3B",X"BC",X"CB",X"B0",X"00",
		X"CC",X"B0",X"3C",X"BB",X"CB",X"00",X"00",X"00",X"00",X"0B",X"BB",X"CB",X"C0",X"00",X"00",X"00",
		X"BB",X"BC",X"0C",X"B0",X"00",X"00",X"00",X"BB",X"C0",X"00",X"00",X"00",X"00",X"00",X"CB",X"BC",
		X"00",X"00",X"00",X"00",X"00",X"02",X"BB",X"C0",X"00",X"00",X"00",X"00",X"BC",X"CB",X"B0",X"00",
		X"00",X"00",X"0B",X"BC",X"BB",X"C0",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"BB",X"00",X"00",X"00",X"0C",X"CB",X"CC",X"B0",X"00",X"00",X"3C",X"BB",X"C3",X"BB",
		X"00",X"00",X"3B",X"BB",X"C0",X"CB",X"00",X"0B",X"3B",X"BB",X"C0",X"BB",X"00",X"0C",X"3B",X"BC",
		X"CC",X"BC",X"00",X"00",X"0B",X"BB",X"3B",X"B0",X"00",X"00",X"0C",X"BB",X"0C",X"B0",X"00",X"00",
		X"00",X"BB",X"C0",X"00",X"00",X"00",X"00",X"BB",X"CB",X"00",X"00",X"00",X"00",X"BB",X"CC",X"00",
		X"00",X"00",X"00",X"BB",X"C0",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"BB",
		X"C0",X"00",X"00",X"00",X"0C",X"BB",X"C0",X"00",X"00",X"00",X"CB",X"BC",X"00",X"00",X"00",X"00",
		X"CB",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"BB",X"00",X"00",X"00",X"0C",X"CC",X"3B",
		X"B0",X"00",X"00",X"0C",X"BC",X"3B",X"B0",X"00",X"00",X"0B",X"BC",X"CB",X"C0",X"00",X"00",X"CB",
		X"CB",X"BB",X"30",X"00",X"CC",X"BC",X"BB",X"BC",X"C0",X"0C",X"BB",X"BC",X"BB",X"3C",X"B0",X"0B",
		X"BC",X"00",X"BB",X"0B",X"B0",X"00",X"BB",X"00",X"00",X"0B",X"B0",X"00",X"0B",X"B0",X"00",X"0B",
		X"C0",X"00",X"0B",X"BB",X"00",X"0B",X"B0",X"00",X"BB",X"C0",X"00",X"0B",X"B0",X"0C",X"BC",X"00",
		X"00",X"CB",X"B0",X"00",X"00",X"00",X"0C",X"BB",X"C0",X"00",X"00",X"00",X"0B",X"BC",X"00",X"00",
		X"00",X"00",X"CC",X"BB",X"00",X"00",X"00",X"00",X"0C",X"CB",X"3C",X"BB",X"00",X"00",X"00",X"3C",
		X"BB",X"C3",X"CB",X"B0",X"00",X"00",X"CB",X"BB",X"CB",X"BB",X"B0",X"0B",X"BC",X"3B",X"BB",X"BB",
		X"BC",X"00",X"0B",X"CC",X"3B",X"BB",X"3C",X"00",X"00",X"0B",X"00",X"BB",X"BB",X"C0",X"00",X"00",
		X"00",X"0B",X"BB",X"CB",X"B0",X"00",X"00",X"00",X"BB",X"B0",X"0B",X"B0",X"00",X"00",X"00",X"BB",
		X"00",X"0B",X"BC",X"BB",X"00",X"00",X"BC",X"00",X"0C",X"BB",X"CB",X"00",X"00",X"BB",X"00",X"00",
		X"0C",X"BB",X"00",X"0C",X"BB",X"00",X"00",X"00",X"BB",X"00",X"CB",X"BB",X"00",X"00",X"00",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"BB",X"B0",X"00",X"00",X"00",
		X"CB",X"BB",X"BB",X"00",X"00",X"3C",X"BB",X"C0",X"CC",X"B0",X"00",X"3B",X"BB",X"00",X"0B",X"B0",
		X"00",X"3B",X"BC",X"30",X"BB",X"00",X"0C",X"3B",X"BC",X"3B",X"B0",X"00",X"0C",X"3B",X"BB",X"3B",
		X"BC",X"00",X"00",X"03",X"BB",X"00",X"CC",X"00",X"00",X"00",X"BB",X"C0",X"00",X"00",X"00",X"00",
		X"BB",X"3C",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"CB",X"B0",X"00",X"00",
		X"00",X"00",X"0B",X"BC",X"00",X"00",X"00",X"00",X"0C",X"BB",X"C0",X"00",X"00",X"00",X"0B",X"BB",
		X"00",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",X"00",X"00",X"03",X"CB",X"B0",X"00",X"00",X"00",
		X"03",X"CC",X"BB",X"BB",X"00",X"00",X"00",X"0C",X"BB",X"B3",X"CC",X"B0",X"00",X"BC",X"0B",X"BB",
		X"BC",X"00",X"CB",X"00",X"BB",X"3B",X"BB",X"BB",X"00",X"BB",X"00",X"00",X"0C",X"B3",X"BB",X"0C",
		X"B0",X"00",X"00",X"03",X"3B",X"BB",X"0B",X"B0",X"00",X"00",X"0C",X"BB",X"C0",X"0C",X"BB",X"00",
		X"00",X"0B",X"B3",X"00",X"00",X"00",X"00",X"00",X"0B",X"BB",X"BB",X"BC",X"00",X"00",X"00",X"00",
		X"33",X"0C",X"BB",X"00",X"00",X"00",X"00",X"CB",X"0C",X"BB",X"00",X"00",X"00",X"0C",X"BB",X"0C",
		X"B0",X"00",X"00",X"00",X"0B",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",
		X"00",X"B0",X"0C",X"00",X"B0",X"00",X"00",X"C0",X"3C",X"3C",X"00",X"00",X"00",X"CB",X"BB",X"C3",
		X"00",X"00",X"0C",X"BB",X"BB",X"B3",X"CB",X"00",X"C7",X"5B",X"BC",X"B3",X"00",X"00",X"B8",X"8B",
		X"BC",X"B3",X"00",X"00",X"78",X"87",X"CC",X"B3",X"CB",X"00",X"C7",X"5C",X"CC",X"B3",X"00",X"00",
		X"00",X"00",X"CC",X"B0",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"A0",X"00",X"00",X"00",X"A0",X"00",X"0A",X"AA",X"A0",X"00",
		X"00",X"A0",X"00",X"00",X"99",X"99",X"AA",X"00",X"A0",X"00",X"A9",X"88",X"88",X"9A",X"AA",X"A0",
		X"00",X"09",X"89",X"78",X"89",X"AA",X"A0",X"00",X"09",X"88",X"88",X"9A",X"00",X"00",X"00",X"A9",
		X"99",X"99",X"AA",X"A0",X"00",X"0A",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"0B",X"BC",X"C0",X"00",
		X"00",X"00",X"BB",X"3B",X"CB",X"00",X"00",X"00",X"BB",X"3B",X"BC",X"C0",X"00",X"00",X"BB",X"CC",
		X"BC",X"BC",X"00",X"00",X"0B",X"BB",X"CC",X"CB",X"B0",X"00",X"CC",X"CB",X"BC",X"0C",X"BB",X"00",
		X"CC",X"CB",X"BC",X"00",X"CB",X"00",X"BB",X"3B",X"BC",X"00",X"B0",X"00",X"BB",X"0C",X"CB",X"00",
		X"00",X"00",X"CB",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"BB",X"C0",X"00",X"00",X"BB",X"00",
		X"CB",X"BC",X"00",X"00",X"BB",X"C0",X"0C",X"BB",X"00",X"00",X"CB",X"BC",X"00",X"00",X"00",X"00",
		X"0C",X"BB",X"00",X"00",X"00",X"00",X"00",X"0B",X"BC",X"00",X"00",X"00",X"00",X"00",X"BB",X"3B",
		X"C0",X"00",X"00",X"00",X"0B",X"B3",X"3B",X"C3",X"BC",X"00",X"00",X"0B",X"B3",X"CB",X"BB",X"CB",
		X"0B",X"B0",X"00",X"BB",X"CC",X"BB",X"3B",X"CB",X"B0",X"00",X"0B",X"CB",X"BC",X"30",X"BC",X"C0",
		X"00",X"CB",X"CB",X"BB",X"00",X"00",X"00",X"00",X"BC",X"0C",X"BB",X"B0",X"00",X"00",X"00",X"00",
		X"00",X"CB",X"B0",X"00",X"00",X"00",X"00",X"0C",X"BB",X"C0",X"00",X"00",X"00",X"00",X"CB",X"B2",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"CC",X"B0",X"00",X"00",X"00",X"00",X"CB",X"BC",X"BB",X"00",
		X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",X"00",X"00",X"0B",X"BC",X"00",X"00",X"00",X"00",X"BC",
		X"CB",X"CC",X"00",X"00",X"0B",X"B3",X"CB",X"BC",X"30",X"00",X"0B",X"C0",X"CB",X"BB",X"30",X"00",
		X"0B",X"B0",X"CB",X"BB",X"3B",X"00",X"0C",X"BC",X"CC",X"BB",X"3C",X"00",X"00",X"BB",X"3B",X"BB",
		X"00",X"00",X"00",X"BC",X"0B",X"BC",X"00",X"00",X"00",X"00",X"CB",X"B0",X"00",X"00",X"00",X"0B",
		X"CB",X"B0",X"00",X"00",X"00",X"0C",X"CB",X"B0",X"00",X"00",X"00",X"00",X"CB",X"B0",X"00",X"00",
		X"00",X"00",X"0B",X"B0",X"00",X"00",X"00",X"00",X"CB",X"B0",X"00",X"00",X"00",X"00",X"CB",X"BC",
		X"00",X"00",X"00",X"00",X"0C",X"BB",X"C0",X"00",X"00",X"00",X"00",X"CB",X"C0",X"00",X"0B",X"BC",
		X"C0",X"00",X"00",X"00",X"BB",X"3C",X"CC",X"00",X"00",X"00",X"BB",X"3C",X"BC",X"00",X"00",X"00",
		X"CB",X"CC",X"BB",X"00",X"00",X"00",X"3B",X"BB",X"CB",X"C0",X"00",X"00",X"CC",X"BB",X"BC",X"BC",
		X"C0",X"00",X"BC",X"3B",X"BC",X"BB",X"BC",X"00",X"BB",X"0B",X"B0",X"0C",X"BB",X"00",X"BB",X"00",
		X"00",X"0B",X"B0",X"00",X"CB",X"00",X"00",X"BB",X"00",X"00",X"BB",X"00",X"0B",X"BB",X"00",X"00",
		X"BB",X"00",X"00",X"CB",X"B0",X"00",X"BB",X"C0",X"00",X"0C",X"BC",X"00",X"CB",X"BC",X"00",X"00",
		X"00",X"00",X"0C",X"BB",X"00",X"00",X"00",X"00",X"00",X"0B",X"BC",X"C0",X"00",X"00",X"00",X"0B",
		X"BC",X"3B",X"CC",X"00",X"00",X"00",X"BB",X"C3",X"CB",X"BC",X"30",X"00",X"00",X"BB",X"BB",X"CB",
		X"BB",X"C0",X"00",X"00",X"0C",X"BB",X"BB",X"BB",X"3C",X"BB",X"00",X"00",X"0C",X"3B",X"BB",X"3C",
		X"CB",X"00",X"00",X"00",X"CB",X"BB",X"B0",X"0B",X"00",X"00",X"00",X"BB",X"CB",X"BB",X"00",X"00",
		X"00",X"00",X"BB",X"00",X"BB",X"B0",X"00",X"0B",X"BC",X"BB",X"00",X"0B",X"B0",X"00",X"0B",X"CB",
		X"BC",X"00",X"0C",X"B0",X"00",X"0B",X"BC",X"00",X"00",X"0B",X"B0",X"00",X"0B",X"B0",X"00",X"00",
		X"0B",X"BC",X"00",X"00",X"00",X"00",X"00",X"0B",X"BB",X"C0",X"00",X"00",X"00",X"00",X"00",X"BB",
		X"B0",X"00",X"BB",X"BC",X"00",X"00",X"00",X"0B",X"BB",X"BB",X"C0",X"00",X"00",X"BC",X"C0",X"CB",
		X"BC",X"30",X"00",X"BB",X"00",X"0B",X"BB",X"30",X"00",X"0B",X"B0",X"3C",X"BB",X"30",X"00",X"00",
		X"BB",X"3C",X"BB",X"3C",X"00",X"0C",X"BB",X"3B",X"BB",X"3C",X"00",X"0C",X"C0",X"0B",X"B3",X"00",
		X"00",X"00",X"00",X"CB",X"B0",X"00",X"00",X"00",X"0C",X"3B",X"B0",X"00",X"00",X"00",X"00",X"0B",
		X"B0",X"00",X"00",X"00",X"00",X"BB",X"C0",X"00",X"00",X"00",X"0C",X"BB",X"00",X"00",X"00",X"00",
		X"CB",X"BC",X"00",X"00",X"00",X"00",X"0B",X"BB",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"00",X"00",X"BB",X"C3",X"00",X"00",X"00",X"00",X"0B",X"BB",X"BC",X"C3",X"00",X"00",X"00",
		X"BC",X"C3",X"BB",X"BC",X"00",X"00",X"0B",X"C0",X"0C",X"BB",X"BB",X"0C",X"B0",X"0B",X"B0",X"0B",
		X"BB",X"BB",X"3B",X"B0",X"00",X"BC",X"0B",X"B3",X"BC",X"00",X"00",X"00",X"BB",X"0B",X"BB",X"33",
		X"00",X"00",X"0B",X"BC",X"00",X"CB",X"BC",X"00",X"00",X"00",X"00",X"00",X"03",X"BB",X"00",X"00",
		X"00",X"0C",X"BB",X"BB",X"BB",X"00",X"00",X"00",X"0B",X"BC",X"03",X"30",X"00",X"00",X"00",X"0B",
		X"BC",X"0B",X"C0",X"00",X"00",X"00",X"00",X"BC",X"0B",X"BC",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"BB",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"B0",X"0C",X"00",X"B0",X"00",X"00",
		X"0C",X"3C",X"30",X"C0",X"00",X"00",X"03",X"CB",X"BB",X"C0",X"00",X"0B",X"C3",X"BB",X"BB",X"BC",
		X"00",X"00",X"03",X"BC",X"BB",X"57",X"C0",X"00",X"03",X"BC",X"BB",X"88",X"B0",X"0B",X"C3",X"BC",
		X"C7",X"88",X"70",X"00",X"03",X"BC",X"CC",X"57",X"C0",X"00",X"00",X"BC",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"A0",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"A0",X"00",X"00",X"AA",X"AA",X"00",X"00",X"A0",X"0A",X"A9",X"99",X"90",
		X"00",X"00",X"AA",X"AA",X"98",X"88",X"89",X"A0",X"00",X"AA",X"A9",X"88",X"79",X"89",X"00",X"00",
		X"00",X"0A",X"98",X"88",X"89",X"00",X"00",X"00",X"AA",X"A9",X"99",X"99",X"A0",X"00",X"00",X"00",
		X"0A",X"AA",X"AA",X"AA",X"00",X"00",X"B0",X"00",X"0C",X"BC",X"00",X"BB",X"BB",X"B0",X"0C",X"BC",
		X"00",X"00",X"B0",X"00",X"00",X"C0",X"00",X"0B",X"CB",X"00",X"CC",X"CC",X"C0",X"0B",X"CB",X"00",
		X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"0B",X"BB",X"BC",X"BB",X"00",X"00",
		X"BB",X"BC",X"BB",X"CC",X"B0",X"00",X"BB",X"3C",X"BC",X"0C",X"C0",X"00",X"BB",X"CC",X"BC",X"3C",
		X"00",X"CB",X"B0",X"CB",X"BB",X"C0",X"00",X"BB",X"0C",X"BB",X"BC",X"C0",X"00",X"BB",X"0B",X"BC",
		X"0C",X"C0",X"00",X"0C",X"0B",X"B0",X"0C",X"B0",X"00",X"00",X"0B",X"B0",X"0B",X"B0",X"00",X"00",
		X"0B",X"B0",X"BB",X"B0",X"00",X"0B",X"CB",X"B0",X"BB",X"B0",X"00",X"0B",X"BB",X"B0",X"0B",X"C0",
		X"00",X"00",X"BB",X"B0",X"00",X"00",X"00",X"00",X"0B",X"C0",X"00",X"00",X"00",X"00",X"00",X"3B",
		X"BB",X"BC",X"00",X"00",X"00",X"BB",X"BC",X"BB",X"C0",X"0B",X"B0",X"CB",X"3C",X"B2",X"C0",X"0B",
		X"BB",X"BB",X"CC",X"BC",X"00",X"00",X"CC",X"BC",X"CB",X"B3",X"00",X"00",X"0C",X"3C",X"BB",X"3C",
		X"00",X"00",X"0B",X"C0",X"00",X"CB",X"00",X"00",X"0B",X"BC",X"00",X"0B",X"00",X"00",X"CB",X"3B",
		X"00",X"0B",X"C0",X"00",X"B3",X"C0",X"00",X"BC",X"B0",X"00",X"BC",X"00",X"00",X"BB",X"B0",X"00",
		X"00",X"00",X"00",X"0B",X"C0",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"0B",X"BB",
		X"B0",X"BB",X"00",X"00",X"00",X"0B",X"BC",X"C0",X"BC",X"00",X"00",X"00",X"0B",X"BC",X"BB",X"2C",
		X"00",X"00",X"00",X"CB",X"BC",X"BB",X"C0",X"00",X"00",X"0B",X"BB",X"BC",X"BB",X"00",X"00",X"00",
		X"BC",X"BC",X"CB",X"CC",X"00",X"00",X"00",X"BC",X"CC",X"C3",X"CC",X"00",X"00",X"00",X"BC",X"00",
		X"0C",X"BB",X"00",X"00",X"BC",X"CB",X"00",X"00",X"CB",X"BB",X"B0",X"CB",X"BB",X"00",X"00",X"00",
		X"CB",X"C0",X"0C",X"BB",X"00",X"00",X"00",X"CB",X"30",X"00",X"BC",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"3B",X"BB",X"B0",X"BB",X"00",X"00",X"00",X"BB",
		X"BC",X"BB",X"CC",X"CC",X"00",X"00",X"BB",X"3C",X"B2",X"00",X"CC",X"00",X"B0",X"BB",X"CC",X"BC",
		X"00",X"BC",X"00",X"BB",X"BC",X"CB",X"BB",X"00",X"CB",X"00",X"CB",X"8C",X"BB",X"B0",X"00",X"00",
		X"00",X"00",X"CB",X"B8",X"CB",X"B0",X"00",X"00",X"00",X"0B",X"B3",X"B3",X"B0",X"00",X"00",X"00",
		X"0B",X"C0",X"B3",X"B0",X"00",X"00",X"00",X"0B",X"B0",X"BB",X"00",X"00",X"00",X"0B",X"CB",X"B0",
		X"00",X"00",X"00",X"00",X"0B",X"BB",X"B0",X"00",X"00",X"00",X"00",X"00",X"BB",X"B0",X"00",X"00",
		X"00",X"00",X"00",X"0B",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"0B",X"BB",X"B0",X"BB",X"00",X"00",X"00",X"BB",X"BC",X"BB",X"CC",X"00",X"00",X"00",
		X"BB",X"3C",X"B2",X"0C",X"00",X"0B",X"B0",X"BB",X"CC",X"B0",X"CC",X"00",X"0B",X"BB",X"BC",X"CB",
		X"B0",X"BC",X"00",X"0C",X"0C",X"CB",X"BB",X"C0",X"00",X"00",X"00",X"0B",X"BB",X"8C",X"C0",X"00",
		X"00",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"0B",X"B0",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"BB",X"BC",X"00",X"00",X"00",X"00",X"00",X"0B",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B3",X"00",X"00",X"00",X"00",X"00",X"0C",X"B3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"0B",X"CB",X"B0",X"BB",X"00",X"00",X"00",X"BB",X"BC",X"BB",X"CB",X"C0",
		X"00",X"00",X"CB",X"BB",X"CC",X"0B",X"C0",X"00",X"00",X"0C",X"BB",X"C0",X"0C",X"C0",X"00",X"0B",
		X"BB",X"BB",X"C3",X"CC",X"00",X"00",X"BB",X"BC",X"CC",X"CB",X"00",X"00",X"00",X"CC",X"CB",X"BB",
		X"CC",X"00",X"00",X"00",X"BB",X"BB",X"B3",X"CC",X"00",X"00",X"00",X"BB",X"00",X"0C",X"B0",X"00",
		X"00",X"00",X"CB",X"00",X"0B",X"B0",X"00",X"00",X"0B",X"BB",X"00",X"0C",X"BB",X"C0",X"00",X"0C",
		X"BB",X"00",X"00",X"B3",X"C0",X"00",X"00",X"00",X"00",X"00",X"B3",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"3B",
		X"BB",X"B0",X"CB",X"00",X"00",X"00",X"0B",X"BB",X"CB",X"CC",X"CB",X"C0",X"00",X"00",X"BB",X"BB",
		X"3B",X"C0",X"0C",X"C0",X"CB",X"BB",X"BB",X"C3",X"CB",X"00",X"0B",X"C0",X"BB",X"B0",X"00",X"CC",
		X"BB",X"C0",X"CB",X"00",X"B0",X"00",X"00",X"CB",X"BB",X"B0",X"CC",X"00",X"00",X"00",X"00",X"0C",
		X"BB",X"00",X"0C",X"00",X"00",X"00",X"00",X"BC",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"BB",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"CB",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"BB",X"C0",X"00",X"00",X"00",X"00",X"00",X"0B",X"B3",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"3C",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"0B",X"00",X"C0",X"0B",X"00",X"00",X"C3",
		X"33",X"C0",X"00",X"5B",X"BB",X"C3",X"30",X"00",X"8B",X"BB",X"BC",X"3C",X"B0",X"77",X"BC",X"BC",
		X"33",X"00",X"5B",X"BC",X"BC",X"30",X"00",X"0B",X"CC",X"BC",X"CC",X"B0",X"00",X"0C",X"BC",X"30",
		X"00",X"00",X"0C",X"BC",X"30",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"0A",X"00",X"00",X"00",
		X"00",X"0A",X"A0",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"0A",X"A0",X"00",X"00",
		X"08",X"9A",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"78",X"9A",X"AA",X"AA",X"A0",X"00",X"00",X"00",
		X"89",X"9A",X"AA",X"A0",X"00",X"00",X"00",X"A9",X"99",X"AA",X"AA",X"AA",X"00",X"00",X"0A",X"AA",
		X"AA",X"AA",X"A0",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"0B",X"BC",X"BB",X"BB",
		X"00",X"00",X"BC",X"CB",X"BC",X"BB",X"B0",X"00",X"CC",X"0C",X"BC",X"3B",X"B0",X"00",X"0C",X"3C",
		X"BC",X"CB",X"B0",X"00",X"00",X"CB",X"BB",X"C0",X"BB",X"C0",X"00",X"CC",X"BB",X"BC",X"0B",X"B0",
		X"00",X"CC",X"0C",X"BB",X"0B",X"B0",X"00",X"BC",X"00",X"BB",X"0C",X"00",X"00",X"BB",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"B0",X"BB",X"00",X"00",X"00",X"BB",X"B0",X"BB",X"CB",X"00",X"00",X"CB",
		X"00",X"BB",X"BB",X"00",X"00",X"00",X"00",X"BB",X"B0",X"00",X"00",X"00",X"00",X"CB",X"00",X"00",
		X"0C",X"BB",X"BB",X"30",X"00",X"00",X"CB",X"BC",X"BB",X"B0",X"00",X"00",X"C2",X"BC",X"3B",X"C0",
		X"BB",X"00",X"0C",X"BC",X"CB",X"BB",X"BB",X"00",X"03",X"BB",X"CC",X"BC",X"C0",X"00",X"0C",X"3B",
		X"BC",X"3C",X"00",X"00",X"0B",X"C0",X"00",X"CB",X"00",X"00",X"0B",X"00",X"0C",X"BB",X"00",X"00",
		X"CB",X"00",X"0B",X"3B",X"C0",X"00",X"BC",X"B0",X"00",X"C3",X"B0",X"00",X"BB",X"B0",X"00",X"0C",
		X"B0",X"00",X"CB",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"0B",
		X"B0",X"BB",X"BB",X"00",X"00",X"00",X"0C",X"B0",X"CC",X"BB",X"00",X"00",X"00",X"0C",X"2B",X"BC",
		X"BB",X"00",X"00",X"00",X"00",X"CB",X"BC",X"BB",X"C0",X"00",X"00",X"00",X"0B",X"BC",X"BB",X"BB",
		X"00",X"00",X"00",X"0C",X"CB",X"CC",X"BC",X"B0",X"00",X"00",X"0C",X"C3",X"CC",X"CC",X"B0",X"00",
		X"00",X"0B",X"BC",X"00",X"0C",X"B0",X"00",X"BB",X"BB",X"C0",X"00",X"0B",X"CC",X"B0",X"CB",X"C0",
		X"00",X"00",X"0B",X"BB",X"C0",X"3B",X"C0",X"00",X"00",X"0B",X"BC",X"00",X"0B",X"B0",X"00",X"00",
		X"0C",X"B0",X"00",X"00",X"0C",X"B0",X"00",X"00",X"00",X"00",X"00",X"0B",X"B0",X"BB",X"BB",X"30",
		X"00",X"0C",X"CC",X"CB",X"BC",X"BB",X"B0",X"00",X"0C",X"C0",X"02",X"BC",X"3B",X"B0",X"00",X"0C",
		X"B0",X"0C",X"BC",X"CB",X"B0",X"B0",X"0B",X"C0",X"0B",X"BB",X"CC",X"BB",X"B0",X"00",X"00",X"00",
		X"BB",X"BC",X"8B",X"C0",X"00",X"00",X"BB",X"C8",X"BB",X"C0",X"00",X"00",X"00",X"B3",X"B3",X"BB",
		X"00",X"00",X"00",X"00",X"B3",X"B0",X"CB",X"00",X"00",X"00",X"00",X"0B",X"B0",X"BB",X"00",X"00",
		X"00",X"00",X"00",X"00",X"BB",X"CB",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",
		X"00",X"00",X"BB",X"B0",X"00",X"00",X"00",X"00",X"00",X"CB",X"00",X"00",X"00",X"B0",X"00",X"00",
		X"00",X"00",X"00",X"0B",X"B0",X"BB",X"BB",X"00",X"00",X"00",X"0C",X"CB",X"BC",X"BB",X"B0",X"00",
		X"00",X"0C",X"02",X"BC",X"3B",X"B0",X"00",X"00",X"0C",X"C0",X"BC",X"CB",X"B0",X"BB",X"00",X"0C",
		X"B0",X"BB",X"CC",X"BB",X"BB",X"00",X"00",X"00",X"CB",X"BB",X"CC",X"0C",X"00",X"00",X"00",X"CC",
		X"8B",X"BB",X"00",X"00",X"00",X"00",X"0C",X"C0",X"0B",X"B0",X"00",X"00",X"00",X"0C",X"C0",X"BB",
		X"00",X"00",X"00",X"00",X"0C",X"BB",X"B0",X"00",X"00",X"00",X"00",X"0B",X"BB",X"00",X"00",X"00",
		X"00",X"00",X"03",X"B0",X"00",X"00",X"00",X"00",X"00",X"03",X"BC",X"00",X"00",X"00",X"00",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"B0",X"BB",X"CB",X"00",X"00",X"00",X"CB",X"CB",X"BC",X"BB",
		X"B0",X"00",X"00",X"CB",X"0C",X"CB",X"BB",X"C0",X"00",X"00",X"CC",X"00",X"CB",X"BC",X"00",X"00",
		X"00",X"0C",X"C3",X"CB",X"BB",X"BB",X"00",X"00",X"00",X"0B",X"CC",X"CC",X"BB",X"B0",X"00",X"00",
		X"0C",X"CB",X"BB",X"CC",X"C0",X"00",X"00",X"0C",X"C3",X"BB",X"BB",X"B0",X"00",X"00",X"00",X"BC",
		X"00",X"0B",X"B0",X"00",X"00",X"00",X"BB",X"00",X"0B",X"C0",X"00",X"00",X"CB",X"BC",X"00",X"0B",
		X"BB",X"00",X"00",X"C3",X"B0",X"00",X"0B",X"BC",X"00",X"00",X"C3",X"B0",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"B0",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",
		X"C0",X"BB",X"BB",X"30",X"00",X"00",X"00",X"CB",X"CC",X"CB",X"CB",X"BB",X"00",X"00",X"00",X"CC",
		X"00",X"CB",X"3B",X"BB",X"B0",X"00",X"00",X"CB",X"00",X"0B",X"C3",X"CB",X"BB",X"BB",X"C0",X"0B",
		X"C0",X"CB",X"BC",X"C0",X"00",X"BB",X"B0",X"0C",X"C0",X"BB",X"BB",X"C0",X"00",X"00",X"B0",X"0C",
		X"00",X"0B",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"BC",X"B0",X"00",X"00",X"00",X"00",
		X"00",X"CB",X"BC",X"C0",X"00",X"00",X"00",X"00",X"0C",X"BB",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"CB",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"3B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"0B",X"00",X"C0",X"0B",
		X"00",X"00",X"C3",X"33",X"C0",X"00",X"00",X"33",X"CB",X"BB",X"50",X"BC",X"3C",X"BB",X"BB",X"80",
		X"03",X"3C",X"BC",X"B7",X"70",X"00",X"3C",X"BC",X"BB",X"50",X"BC",X"CC",X"BC",X"CB",X"00",X"00",
		X"3C",X"BC",X"00",X"00",X"00",X"3C",X"BC",X"00",X"00",X"0A",X"00",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"0A",X"A0",X"00",X"00",
		X"00",X"0A",X"AA",X"AA",X"AA",X"98",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"98",X"70",X"00",
		X"00",X"00",X"00",X"AA",X"AA",X"99",X"80",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"A9",X"99",X"A0",
		X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"90",X"00",X"0A",X"9A",X"00",X"99",
		X"99",X"90",X"0A",X"9A",X"00",X"00",X"90",X"00",X"00",X"A0",X"00",X"09",X"A9",X"00",X"AA",X"AA",
		X"A0",X"09",X"A9",X"00",X"00",X"A0",X"00",X"09",X"9A",X"A0",X"00",X"00",X"00",X"99",X"39",X"A9",
		X"00",X"00",X"00",X"99",X"39",X"9A",X"A0",X"00",X"00",X"99",X"AA",X"9A",X"9A",X"00",X"00",X"09",
		X"99",X"AA",X"A9",X"90",X"00",X"AA",X"A9",X"9A",X"0A",X"99",X"00",X"AA",X"A9",X"9A",X"00",X"A9",
		X"00",X"99",X"39",X"9A",X"00",X"90",X"00",X"99",X"0A",X"A9",X"00",X"00",X"00",X"A9",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"99",X"A0",X"00",X"00",X"99",X"00",X"A9",X"9A",X"00",X"00",X"99",
		X"A0",X"0A",X"99",X"00",X"00",X"A9",X"9A",X"00",X"00",X"00",X"00",X"0A",X"99",X"00",X"00",X"00",
		X"00",X"00",X"09",X"9A",X"00",X"00",X"00",X"00",X"00",X"99",X"39",X"A0",X"00",X"00",X"00",X"09",
		X"93",X"39",X"A3",X"9A",X"00",X"00",X"09",X"93",X"A9",X"99",X"A9",X"09",X"90",X"00",X"99",X"AA",
		X"99",X"39",X"A9",X"90",X"00",X"09",X"A9",X"9A",X"30",X"9A",X"A0",X"00",X"A9",X"A9",X"99",X"00",
		X"00",X"00",X"00",X"9A",X"0A",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"A9",X"90",X"00",X"00",
		X"00",X"00",X"0A",X"99",X"A0",X"00",X"00",X"00",X"00",X"A9",X"92",X"00",X"00",X"00",X"00",X"00",
		X"99",X"AA",X"90",X"00",X"00",X"00",X"00",X"A9",X"9A",X"99",X"00",X"00",X"00",X"00",X"09",X"90",
		X"00",X"00",X"00",X"00",X"09",X"9A",X"00",X"00",X"00",X"00",X"9A",X"A9",X"AA",X"00",X"00",X"09",
		X"93",X"A9",X"9A",X"30",X"00",X"09",X"A0",X"A9",X"99",X"30",X"00",X"09",X"90",X"A9",X"99",X"39",
		X"00",X"0A",X"9A",X"AA",X"99",X"3A",X"00",X"00",X"99",X"39",X"99",X"00",X"00",X"00",X"9A",X"09",
		X"9A",X"00",X"00",X"00",X"00",X"A9",X"90",X"00",X"00",X"00",X"09",X"A9",X"90",X"00",X"00",X"00",
		X"0A",X"A9",X"90",X"00",X"00",X"00",X"00",X"A9",X"90",X"00",X"00",X"00",X"00",X"09",X"90",X"00",
		X"00",X"00",X"00",X"A9",X"90",X"00",X"00",X"00",X"00",X"A9",X"9A",X"00",X"00",X"00",X"00",X"0A",
		X"99",X"A0",X"00",X"00",X"00",X"00",X"A9",X"A0",X"00",X"09",X"9A",X"A0",X"00",X"00",X"00",X"99",
		X"3A",X"AA",X"00",X"00",X"00",X"99",X"3A",X"9A",X"00",X"00",X"00",X"A9",X"AA",X"99",X"00",X"00",
		X"00",X"39",X"99",X"A9",X"A0",X"00",X"00",X"AA",X"99",X"9A",X"9A",X"A0",X"00",X"9A",X"39",X"9A",
		X"99",X"9A",X"00",X"99",X"09",X"90",X"0A",X"99",X"00",X"99",X"00",X"00",X"09",X"90",X"00",X"A9",
		X"00",X"00",X"99",X"00",X"00",X"99",X"00",X"09",X"99",X"00",X"00",X"99",X"00",X"00",X"A9",X"90",
		X"00",X"99",X"A0",X"00",X"0A",X"9A",X"00",X"A9",X"9A",X"00",X"00",X"00",X"00",X"0A",X"99",X"00",
		X"00",X"00",X"00",X"00",X"09",X"9A",X"A0",X"00",X"00",X"00",X"09",X"9A",X"39",X"AA",X"00",X"00",
		X"00",X"99",X"A3",X"A9",X"9A",X"30",X"00",X"00",X"99",X"99",X"A9",X"99",X"A0",X"00",X"00",X"0A",
		X"99",X"99",X"99",X"3A",X"99",X"00",X"00",X"0A",X"39",X"99",X"3A",X"A9",X"00",X"00",X"00",X"A9",
		X"99",X"90",X"09",X"00",X"00",X"00",X"99",X"A9",X"99",X"00",X"00",X"00",X"00",X"99",X"00",X"99",
		X"90",X"00",X"09",X"9A",X"99",X"00",X"09",X"90",X"00",X"09",X"A9",X"9A",X"00",X"0A",X"90",X"00",
		X"09",X"9A",X"00",X"00",X"09",X"90",X"00",X"09",X"90",X"00",X"00",X"09",X"9A",X"00",X"00",X"00",
		X"00",X"00",X"09",X"99",X"A0",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"99",X"9A",X"00",
		X"00",X"00",X"09",X"99",X"99",X"A0",X"00",X"00",X"9A",X"A0",X"A9",X"9A",X"30",X"00",X"99",X"00",
		X"09",X"99",X"30",X"00",X"09",X"90",X"3A",X"99",X"30",X"00",X"00",X"99",X"3A",X"99",X"3A",X"00",
		X"0A",X"99",X"39",X"99",X"3A",X"00",X"0A",X"A0",X"09",X"93",X"00",X"00",X"00",X"00",X"A9",X"90",
		X"00",X"00",X"00",X"0A",X"39",X"90",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"00",X"00",X"00",
		X"99",X"A0",X"00",X"00",X"00",X"0A",X"99",X"00",X"00",X"00",X"00",X"A9",X"9A",X"00",X"00",X"00",
		X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"99",X"A3",
		X"00",X"00",X"00",X"00",X"09",X"99",X"9A",X"A3",X"00",X"00",X"00",X"9A",X"A3",X"99",X"9A",X"00",
		X"00",X"09",X"A0",X"0A",X"99",X"99",X"0A",X"90",X"09",X"90",X"09",X"99",X"99",X"39",X"90",X"00",
		X"9A",X"09",X"93",X"9A",X"00",X"00",X"00",X"99",X"09",X"99",X"33",X"00",X"00",X"09",X"9A",X"00",
		X"A9",X"9A",X"00",X"00",X"00",X"00",X"00",X"03",X"99",X"00",X"00",X"00",X"0A",X"99",X"99",X"99",
		X"00",X"00",X"00",X"09",X"9A",X"03",X"30",X"00",X"00",X"00",X"09",X"9A",X"09",X"A0",X"00",X"00",
		X"00",X"00",X"9A",X"09",X"9A",X"00",X"00",X"00",X"00",X"00",X"0A",X"99",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"90",X"0A",X"00",X"90",X"00",X"00",X"0A",X"3A",X"30",X"A0",X"00",
		X"00",X"03",X"A9",X"99",X"A0",X"00",X"09",X"A3",X"99",X"99",X"9A",X"00",X"00",X"03",X"9A",X"99",
		X"57",X"A0",X"00",X"03",X"9A",X"99",X"88",X"90",X"09",X"A3",X"9A",X"A7",X"88",X"70",X"00",X"03",
		X"9A",X"AA",X"57",X"A0",X"00",X"00",X"9A",X"A0",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"09",X"9A",X"99",X"99",X"00",X"00",X"9A",X"A9",X"9A",X"99",X"90",X"00",X"AA",X"0A",X"9A",X"39",
		X"90",X"00",X"0A",X"3A",X"9A",X"A9",X"90",X"00",X"00",X"A9",X"99",X"A0",X"99",X"A0",X"00",X"AA",
		X"99",X"9A",X"09",X"90",X"00",X"AA",X"0A",X"99",X"09",X"90",X"00",X"9A",X"00",X"99",X"0A",X"00",
		X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"99",X"00",X"00",X"00",X"99",X"90",X"99",
		X"A9",X"00",X"00",X"A9",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"00",
		X"00",X"A9",X"00",X"00",X"0A",X"99",X"99",X"30",X"00",X"00",X"A9",X"9A",X"99",X"90",X"00",X"00",
		X"A2",X"9A",X"39",X"A0",X"99",X"00",X"0A",X"9A",X"A9",X"99",X"99",X"00",X"03",X"99",X"AA",X"9A",
		X"A0",X"00",X"0A",X"39",X"9A",X"3A",X"00",X"00",X"09",X"A0",X"00",X"A9",X"00",X"00",X"09",X"00",
		X"0A",X"99",X"00",X"00",X"A9",X"00",X"09",X"39",X"A0",X"00",X"9A",X"90",X"00",X"A3",X"90",X"00",
		X"99",X"90",X"00",X"0A",X"90",X"00",X"A9",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"09",X"90",X"99",X"99",X"00",X"00",X"00",X"0A",X"90",X"AA",X"99",X"00",X"00",
		X"00",X"0A",X"29",X"9A",X"99",X"00",X"00",X"00",X"00",X"A9",X"9A",X"99",X"A0",X"00",X"00",X"00",
		X"09",X"9A",X"99",X"99",X"00",X"00",X"00",X"0A",X"A9",X"AA",X"9A",X"90",X"00",X"00",X"0A",X"A3",
		X"AA",X"AA",X"90",X"00",X"00",X"09",X"9A",X"00",X"0A",X"90",X"00",X"99",X"99",X"A0",X"00",X"09",
		X"AA",X"90",X"A9",X"A0",X"00",X"00",X"09",X"99",X"A0",X"39",X"A0",X"00",X"00",X"09",X"9A",X"00",
		X"09",X"90",X"00",X"00",X"0A",X"90",X"00",X"00",X"0A",X"90",X"00",X"00",X"00",X"00",X"00",X"09",
		X"90",X"99",X"99",X"30",X"00",X"0A",X"AA",X"A9",X"9A",X"99",X"90",X"00",X"0A",X"A0",X"02",X"9A",
		X"39",X"90",X"00",X"0A",X"90",X"0A",X"9A",X"A9",X"90",X"90",X"09",X"A0",X"09",X"99",X"AA",X"99",
		X"90",X"00",X"00",X"00",X"99",X"9A",X"89",X"A0",X"00",X"00",X"99",X"A8",X"99",X"A0",X"00",X"00",
		X"00",X"93",X"93",X"99",X"00",X"00",X"00",X"00",X"93",X"90",X"A9",X"00",X"00",X"00",X"00",X"09",
		X"90",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"A9",X"00",X"00",X"00",X"00",X"00",X"99",
		X"99",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"A9",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"99",X"99",X"00",X"00",X"00",X"0A",X"A9",
		X"9A",X"99",X"90",X"00",X"00",X"0A",X"02",X"9A",X"39",X"90",X"00",X"00",X"0A",X"A0",X"9A",X"A9",
		X"90",X"99",X"00",X"0A",X"90",X"99",X"AA",X"99",X"99",X"00",X"00",X"00",X"A9",X"99",X"AA",X"0A",
		X"00",X"00",X"00",X"AA",X"89",X"99",X"00",X"00",X"00",X"00",X"0A",X"A0",X"09",X"90",X"00",X"00",
		X"00",X"0A",X"A0",X"99",X"00",X"00",X"00",X"00",X"0A",X"99",X"90",X"00",X"00",X"00",X"00",X"09",
		X"99",X"00",X"00",X"00",X"00",X"00",X"03",X"90",X"00",X"00",X"00",X"00",X"00",X"03",X"9A",X"00",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"99",X"A9",X"00",X"00",X"00",
		X"A9",X"A9",X"9A",X"99",X"90",X"00",X"00",X"A9",X"0A",X"A9",X"99",X"A0",X"00",X"00",X"AA",X"00",
		X"A9",X"9A",X"00",X"00",X"00",X"0A",X"A3",X"A9",X"99",X"99",X"00",X"00",X"00",X"09",X"AA",X"AA",
		X"99",X"90",X"00",X"00",X"0A",X"A9",X"99",X"AA",X"A0",X"00",X"00",X"0A",X"A3",X"99",X"99",X"90",
		X"00",X"00",X"00",X"9A",X"00",X"09",X"90",X"00",X"00",X"00",X"99",X"00",X"09",X"A0",X"00",X"00",
		X"A9",X"9A",X"00",X"09",X"99",X"00",X"00",X"A3",X"90",X"00",X"09",X"9A",X"00",X"00",X"A3",X"90",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"90",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"A0",X"99",X"99",X"30",X"00",X"00",X"00",X"A9",X"AA",X"A9",X"A9",X"99",
		X"00",X"00",X"00",X"AA",X"00",X"A9",X"39",X"99",X"90",X"00",X"00",X"A9",X"00",X"09",X"A3",X"A9",
		X"99",X"99",X"A0",X"09",X"A0",X"A9",X"9A",X"A0",X"00",X"99",X"90",X"0A",X"A0",X"99",X"99",X"A0",
		X"00",X"00",X"90",X"0A",X"00",X"09",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"9A",X"90",
		X"00",X"00",X"00",X"00",X"00",X"A9",X"9A",X"A0",X"00",X"00",X"00",X"00",X"0A",X"99",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"A9",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"A3",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"09",X"00",X"A0",X"09",X"00",X"00",X"A3",X"33",X"A0",X"00",X"00",X"33",X"A9",X"99",X"50",X"9A",
		X"3A",X"99",X"99",X"80",X"03",X"3A",X"9A",X"97",X"70",X"00",X"3A",X"9A",X"99",X"50",X"9A",X"AA",
		X"9A",X"A9",X"00",X"00",X"3A",X"9A",X"00",X"00",X"00",X"3A",X"9A",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"99",X"00",X"00",X"00",X"09",X"A9",X"39",X"90",X"00",X"00",X"AA",X"99",X"39",X"90",X"00",
		X"0A",X"9A",X"9A",X"A9",X"90",X"00",X"99",X"AA",X"A9",X"99",X"00",X"09",X"9A",X"0A",X"99",X"AA",
		X"A0",X"09",X"A0",X"0A",X"99",X"AA",X"A0",X"00",X"90",X"0A",X"99",X"39",X"90",X"00",X"00",X"09",
		X"AA",X"09",X"90",X"00",X"00",X"09",X"90",X"09",X"A0",X"00",X"00",X"A9",X"90",X"09",X"90",X"00",
		X"0A",X"99",X"A0",X"09",X"90",X"00",X"09",X"9A",X"00",X"A9",X"90",X"00",X"00",X"00",X"0A",X"99",
		X"A0",X"00",X"00",X"00",X"09",X"9A",X"00",X"00",X"00",X"00",X"0A",X"99",X"00",X"00",X"00",X"00",
		X"00",X"A9",X"39",X"90",X"00",X"00",X"0A",X"93",X"A9",X"33",X"99",X"00",X"99",X"09",X"A9",X"99",
		X"A3",X"99",X"00",X"99",X"A9",X"39",X"9A",X"A9",X"90",X"00",X"AA",X"90",X"3A",X"99",X"A9",X"00",
		X"00",X"00",X"00",X"09",X"99",X"A9",X"A0",X"00",X"00",X"00",X"99",X"9A",X"0A",X"90",X"00",X"00",
		X"00",X"99",X"A0",X"00",X"00",X"00",X"00",X"00",X"A9",X"9A",X"00",X"00",X"00",X"00",X"00",X"02",
		X"99",X"A0",X"00",X"00",X"00",X"00",X"9A",X"A9",X"90",X"00",X"00",X"00",X"09",X"9A",X"99",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"0A",X"99",X"00",X"00",X"00",
		X"0A",X"A9",X"AA",X"90",X"00",X"00",X"3A",X"99",X"A3",X"99",X"00",X"00",X"39",X"99",X"A0",X"A9",
		X"00",X"09",X"39",X"99",X"A0",X"99",X"00",X"0A",X"39",X"9A",X"AA",X"9A",X"00",X"00",X"09",X"99",
		X"39",X"90",X"00",X"00",X"0A",X"99",X"0A",X"90",X"00",X"00",X"00",X"99",X"A0",X"00",X"00",X"00",
		X"00",X"99",X"A9",X"00",X"00",X"00",X"00",X"99",X"AA",X"00",X"00",X"00",X"00",X"99",X"A0",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"99",X"A0",X"00",X"00",X"00",X"0A",X"99",
		X"A0",X"00",X"00",X"00",X"A9",X"9A",X"00",X"00",X"00",X"00",X"A9",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"99",X"00",X"00",X"00",X"0A",X"AA",X"39",X"90",X"00",X"00",X"0A",X"9A",X"39",
		X"90",X"00",X"00",X"09",X"9A",X"A9",X"A0",X"00",X"00",X"A9",X"A9",X"99",X"30",X"00",X"AA",X"9A",
		X"99",X"9A",X"A0",X"0A",X"99",X"9A",X"99",X"3A",X"90",X"09",X"9A",X"00",X"99",X"09",X"90",X"00",
		X"99",X"00",X"00",X"09",X"90",X"00",X"09",X"90",X"00",X"09",X"A0",X"00",X"09",X"99",X"00",X"09",
		X"90",X"00",X"99",X"A0",X"00",X"09",X"90",X"0A",X"9A",X"00",X"00",X"A9",X"90",X"00",X"00",X"00",
		X"0A",X"99",X"A0",X"00",X"00",X"00",X"09",X"9A",X"00",X"00",X"00",X"00",X"AA",X"99",X"00",X"00",
		X"00",X"00",X"0A",X"A9",X"3A",X"99",X"00",X"00",X"00",X"3A",X"99",X"A3",X"A9",X"90",X"00",X"00",
		X"A9",X"99",X"A9",X"99",X"90",X"09",X"9A",X"39",X"99",X"99",X"9A",X"00",X"09",X"AA",X"39",X"99",
		X"3A",X"00",X"00",X"09",X"00",X"99",X"99",X"A0",X"00",X"00",X"00",X"09",X"99",X"A9",X"90",X"00",
		X"00",X"00",X"99",X"90",X"09",X"90",X"00",X"00",X"00",X"99",X"00",X"09",X"9A",X"99",X"00",X"00",
		X"9A",X"00",X"0A",X"99",X"A9",X"00",X"00",X"99",X"00",X"00",X"0A",X"99",X"00",X"0A",X"99",X"00",
		X"00",X"00",X"99",X"00",X"A9",X"99",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"99",X"90",X"00",X"00",X"00",X"A9",X"99",X"99",X"00",X"00",X"3A",
		X"99",X"A0",X"AA",X"90",X"00",X"39",X"99",X"00",X"09",X"90",X"00",X"39",X"9A",X"30",X"99",X"00",
		X"0A",X"39",X"9A",X"39",X"90",X"00",X"0A",X"39",X"99",X"39",X"9A",X"00",X"00",X"03",X"99",X"00",
		X"AA",X"00",X"00",X"00",X"99",X"A0",X"00",X"00",X"00",X"00",X"99",X"3A",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"00",X"00",X"A9",X"90",X"00",X"00",X"00",X"00",X"09",X"9A",X"00",X"00",
		X"00",X"00",X"0A",X"99",X"A0",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"09",X"90",
		X"00",X"00",X"00",X"00",X"03",X"A9",X"90",X"00",X"00",X"00",X"03",X"AA",X"99",X"99",X"00",X"00",
		X"00",X"0A",X"99",X"93",X"AA",X"90",X"00",X"9A",X"09",X"99",X"9A",X"00",X"A9",X"00",X"99",X"39",
		X"99",X"99",X"00",X"99",X"00",X"00",X"0A",X"93",X"99",X"0A",X"90",X"00",X"00",X"03",X"39",X"99",
		X"09",X"90",X"00",X"00",X"0A",X"99",X"A0",X"0A",X"99",X"00",X"00",X"09",X"93",X"00",X"00",X"00",
		X"00",X"00",X"09",X"99",X"99",X"9A",X"00",X"00",X"00",X"00",X"33",X"0A",X"99",X"00",X"00",X"00",
		X"00",X"A9",X"0A",X"99",X"00",X"00",X"00",X"0A",X"99",X"0A",X"90",X"00",X"00",X"00",X"09",X"9A",
		X"00",X"00",X"00",X"00",X"20",X"49",X"4E",X"46",X"45",X"52",X"4E",X"4F",X"20",X"2D",X"20",X"43",
		X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",X"38",
		X"34",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",
		X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"90",X"0A",X"00",X"90",X"00",X"00",X"A0",X"3A",X"3A",X"00",X"00",X"00",X"A9",X"99",
		X"A3",X"00",X"00",X"0A",X"99",X"99",X"93",X"A9",X"00",X"A7",X"59",X"9A",X"93",X"00",X"00",X"98",
		X"89",X"9A",X"93",X"00",X"00",X"78",X"87",X"AA",X"93",X"A9",X"00",X"A7",X"5A",X"AA",X"93",X"00",
		X"00",X"00",X"00",X"AA",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"99",
		X"9A",X"99",X"00",X"00",X"99",X"9A",X"99",X"AA",X"90",X"00",X"99",X"3A",X"9A",X"0A",X"A0",X"00",
		X"99",X"AA",X"9A",X"3A",X"00",X"A9",X"90",X"A9",X"99",X"A0",X"00",X"99",X"0A",X"99",X"9A",X"A0",
		X"00",X"99",X"09",X"9A",X"0A",X"A0",X"00",X"0A",X"09",X"90",X"0A",X"90",X"00",X"00",X"09",X"90",
		X"09",X"90",X"00",X"00",X"09",X"90",X"99",X"90",X"00",X"09",X"A9",X"90",X"99",X"90",X"00",X"09",
		X"99",X"90",X"09",X"A0",X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"09",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"39",X"99",X"9A",X"00",X"00",X"00",X"99",X"9A",X"99",X"A0",X"09",X"90",X"A9",
		X"3A",X"92",X"A0",X"09",X"99",X"99",X"AA",X"9A",X"00",X"00",X"AA",X"9A",X"A9",X"93",X"00",X"00",
		X"0A",X"3A",X"99",X"3A",X"00",X"00",X"09",X"A0",X"00",X"A9",X"00",X"00",X"09",X"9A",X"00",X"09",
		X"00",X"00",X"A9",X"39",X"00",X"09",X"A0",X"00",X"93",X"A0",X"00",X"9A",X"90",X"00",X"9A",X"00",
		X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"09",X"A0",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"09",X"99",X"90",X"99",X"00",X"00",X"00",X"09",X"9A",X"A0",X"9A",X"00",X"00",X"00",
		X"09",X"9A",X"99",X"2A",X"00",X"00",X"00",X"A9",X"9A",X"99",X"A0",X"00",X"00",X"09",X"99",X"9A",
		X"99",X"00",X"00",X"00",X"9A",X"9A",X"A9",X"AA",X"00",X"00",X"00",X"9A",X"AA",X"A3",X"AA",X"00",
		X"00",X"00",X"9A",X"00",X"0A",X"99",X"00",X"00",X"9A",X"A9",X"00",X"00",X"A9",X"99",X"90",X"A9",
		X"99",X"00",X"00",X"00",X"A9",X"A0",X"0A",X"99",X"00",X"00",X"00",X"A9",X"30",X"00",X"9A",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"39",X"99",X"90",X"99",
		X"00",X"00",X"00",X"99",X"9A",X"99",X"AA",X"AA",X"00",X"00",X"99",X"3A",X"92",X"00",X"AA",X"00",
		X"90",X"99",X"AA",X"9A",X"00",X"9A",X"00",X"99",X"9A",X"A9",X"99",X"00",X"A9",X"00",X"A9",X"8A",
		X"99",X"90",X"00",X"00",X"00",X"00",X"A9",X"98",X"A9",X"90",X"00",X"00",X"00",X"09",X"93",X"93",
		X"90",X"00",X"00",X"00",X"09",X"A0",X"93",X"90",X"00",X"00",X"00",X"09",X"90",X"99",X"00",X"00",
		X"00",X"09",X"A9",X"90",X"00",X"00",X"00",X"00",X"09",X"99",X"90",X"00",X"00",X"00",X"00",X"00",
		X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"99",X"90",X"99",X"00",X"00",X"00",X"99",X"9A",X"99",
		X"AA",X"00",X"00",X"00",X"99",X"3A",X"92",X"0A",X"00",X"09",X"90",X"99",X"AA",X"90",X"AA",X"00",
		X"09",X"99",X"9A",X"A9",X"90",X"9A",X"00",X"0A",X"0A",X"A9",X"99",X"A0",X"00",X"00",X"00",X"09",
		X"99",X"8A",X"A0",X"00",X"00",X"00",X"99",X"00",X"AA",X"00",X"00",X"00",X"00",X"09",X"90",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"99",X"9A",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"00",X"00",X"0A",X"93",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"A9",X"90",X"99",X"00",X"00",X"00",X"99",
		X"9A",X"99",X"A9",X"A0",X"00",X"00",X"A9",X"99",X"AA",X"09",X"A0",X"00",X"00",X"0A",X"99",X"A0",
		X"0A",X"A0",X"00",X"09",X"99",X"99",X"A3",X"AA",X"00",X"00",X"99",X"9A",X"AA",X"A9",X"00",X"00",
		X"00",X"AA",X"A9",X"99",X"AA",X"00",X"00",X"00",X"99",X"99",X"93",X"AA",X"00",X"00",X"00",X"99",
		X"00",X"0A",X"90",X"00",X"00",X"00",X"A9",X"00",X"09",X"90",X"00",X"00",X"09",X"99",X"00",X"0A",
		X"99",X"A0",X"00",X"0A",X"99",X"00",X"00",X"93",X"A0",X"00",X"00",X"00",X"00",X"00",X"93",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"39",X"99",X"90",X"A9",X"00",X"00",X"00",X"09",X"99",X"A9",X"AA",X"A9",X"A0",
		X"00",X"00",X"99",X"99",X"39",X"A0",X"0A",X"A0",X"A9",X"99",X"99",X"A3",X"A9",X"00",X"09",X"A0",
		X"99",X"90",X"00",X"AA",X"99",X"A0",X"A9",X"00",X"90",X"00",X"00",X"A9",X"99",X"90",X"AA",X"00",
		X"00",X"00",X"00",X"0A",X"99",X"00",X"0A",X"00",X"00",X"00",X"00",X"9A",X"9A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"99",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"9A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"99",X"A0",X"00",X"00",X"00",X"00",X"00",X"09",X"93",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"09",X"3A",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"00",X"A0",
		X"09",X"00",X"00",X"A3",X"33",X"A0",X"00",X"59",X"99",X"A3",X"30",X"00",X"89",X"99",X"9A",X"3A",
		X"90",X"77",X"9A",X"9A",X"33",X"00",X"59",X"9A",X"9A",X"30",X"00",X"09",X"AA",X"9A",X"AA",X"90",
		X"00",X"0A",X"9A",X"30",X"00",X"00",X"0A",X"9A",X"30",X"00",X"00",X"E0",X"00",X"0F",X"EF",X"00",
		X"EE",X"EE",X"E0",X"0F",X"EF",X"00",X"00",X"E0",X"00",X"00",X"F0",X"00",X"0E",X"FE",X"00",X"FF",
		X"FF",X"F0",X"0E",X"FE",X"00",X"00",X"F0",X"00",X"0E",X"EF",X"F0",X"00",X"00",X"00",X"EE",X"3E",
		X"FE",X"00",X"00",X"00",X"EE",X"3E",X"EF",X"F0",X"00",X"00",X"EE",X"FF",X"EF",X"EF",X"00",X"00",
		X"0E",X"EE",X"FF",X"FE",X"E0",X"00",X"FF",X"FE",X"EF",X"0F",X"EE",X"00",X"FF",X"FE",X"EF",X"00",
		X"FE",X"00",X"EE",X"3E",X"EF",X"00",X"E0",X"00",X"EE",X"0F",X"FE",X"00",X"00",X"00",X"FE",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"00",X"EE",X"F0",X"00",X"00",X"EE",X"00",X"FE",X"EF",X"00",X"00",
		X"EE",X"F0",X"0F",X"EE",X"00",X"00",X"FE",X"EF",X"00",X"00",X"00",X"00",X"0F",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"EF",X"00",X"00",X"00",X"00",X"00",X"EE",X"3E",X"F0",X"00",X"00",X"00",
		X"0E",X"E3",X"3E",X"F3",X"EF",X"00",X"00",X"0E",X"E3",X"FE",X"EE",X"FE",X"0E",X"E0",X"00",X"EE",
		X"FF",X"EE",X"3E",X"FE",X"E0",X"00",X"0E",X"FE",X"EF",X"30",X"EF",X"F0",X"00",X"FE",X"FE",X"EE",
		X"00",X"00",X"00",X"00",X"EF",X"0F",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"FE",X"E0",X"00",
		X"00",X"00",X"00",X"0F",X"EE",X"F0",X"00",X"00",X"00",X"00",X"FE",X"E2",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"FF",X"E0",X"00",X"00",X"00",X"00",X"FE",X"EF",X"EE",X"00",X"00",X"00",X"00",X"0E",
		X"E0",X"00",X"00",X"00",X"00",X"0E",X"EF",X"00",X"00",X"00",X"00",X"EF",X"FE",X"FF",X"00",X"00",
		X"0E",X"E3",X"FE",X"EF",X"30",X"00",X"0E",X"F0",X"FE",X"EE",X"30",X"00",X"0E",X"E0",X"FE",X"EE",
		X"3E",X"00",X"0F",X"EF",X"FF",X"EE",X"3F",X"00",X"00",X"EE",X"3E",X"EE",X"00",X"00",X"00",X"EF",
		X"0E",X"EF",X"00",X"00",X"00",X"00",X"FE",X"E0",X"00",X"00",X"00",X"0E",X"FE",X"E0",X"00",X"00",
		X"00",X"0F",X"FE",X"E0",X"00",X"00",X"00",X"00",X"FE",X"E0",X"00",X"00",X"00",X"00",X"0E",X"E0",
		X"00",X"00",X"00",X"00",X"FE",X"E0",X"00",X"00",X"00",X"00",X"FE",X"EF",X"00",X"00",X"00",X"00",
		X"0F",X"EE",X"F0",X"00",X"00",X"00",X"00",X"FE",X"F0",X"00",X"0E",X"EF",X"F0",X"00",X"00",X"00",
		X"EE",X"3F",X"FF",X"00",X"00",X"00",X"EE",X"3F",X"EF",X"00",X"00",X"00",X"FE",X"FF",X"EE",X"00",
		X"00",X"00",X"3E",X"EE",X"FE",X"F0",X"00",X"00",X"FF",X"EE",X"EF",X"EF",X"F0",X"00",X"EF",X"3E",
		X"EF",X"EE",X"EF",X"00",X"EE",X"0E",X"E0",X"0F",X"EE",X"00",X"EE",X"00",X"00",X"0E",X"E0",X"00",
		X"FE",X"00",X"00",X"EE",X"00",X"00",X"EE",X"00",X"0E",X"EE",X"00",X"00",X"EE",X"00",X"00",X"FE",
		X"E0",X"00",X"EE",X"F0",X"00",X"0F",X"EF",X"00",X"FE",X"EF",X"00",X"00",X"00",X"00",X"0F",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"EF",X"F0",X"00",X"00",X"00",X"0E",X"EF",X"3E",X"FF",X"00",
		X"00",X"00",X"EE",X"F3",X"FE",X"EF",X"30",X"00",X"00",X"EE",X"EE",X"FE",X"EE",X"F0",X"00",X"00",
		X"0F",X"EE",X"EE",X"EE",X"3F",X"EE",X"00",X"00",X"0F",X"3E",X"EE",X"3F",X"FE",X"00",X"00",X"00",
		X"FE",X"EE",X"E0",X"0E",X"00",X"00",X"00",X"EE",X"FE",X"EE",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"EE",X"E0",X"00",X"0E",X"EF",X"EE",X"00",X"0E",X"E0",X"00",X"0E",X"FE",X"EF",X"00",X"0F",X"E0",
		X"00",X"0E",X"EF",X"00",X"00",X"0E",X"E0",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"EF",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"EE",X"F0",X"00",X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",X"EE",X"EF",
		X"00",X"00",X"00",X"0E",X"EE",X"EE",X"F0",X"00",X"00",X"EF",X"F0",X"FE",X"EF",X"30",X"00",X"EE",
		X"00",X"0E",X"EE",X"30",X"00",X"0E",X"E0",X"3F",X"EE",X"30",X"00",X"00",X"EE",X"3F",X"EE",X"3F",
		X"00",X"0F",X"EE",X"3E",X"EE",X"3F",X"00",X"0F",X"F0",X"0E",X"E3",X"00",X"00",X"00",X"00",X"FE",
		X"E0",X"00",X"00",X"00",X"0F",X"3E",X"E0",X"00",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",
		X"00",X"EE",X"F0",X"00",X"00",X"00",X"0F",X"EE",X"00",X"00",X"00",X"00",X"FE",X"EF",X"00",X"00",
		X"00",X"00",X"0E",X"EE",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"F3",X"00",X"00",X"00",X"00",X"0E",X"EE",X"EF",X"F3",X"00",X"00",X"00",X"EF",X"F3",X"EE",X"EF",
		X"00",X"00",X"0E",X"F0",X"0F",X"EE",X"EE",X"0F",X"E0",X"0E",X"E0",X"0E",X"EE",X"EE",X"3E",X"E0",
		X"00",X"EF",X"0E",X"E3",X"EF",X"00",X"00",X"00",X"EE",X"0E",X"EE",X"33",X"00",X"00",X"0E",X"EF",
		X"00",X"FE",X"EF",X"00",X"00",X"00",X"00",X"00",X"03",X"EE",X"00",X"00",X"00",X"0F",X"EE",X"EE",
		X"EE",X"00",X"00",X"00",X"0E",X"EF",X"03",X"30",X"00",X"00",X"00",X"0E",X"EF",X"0E",X"F0",X"00",
		X"00",X"00",X"00",X"EF",X"0E",X"EF",X"00",X"00",X"00",X"00",X"00",X"0F",X"EE",X"00",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"E0",X"0F",X"00",X"E0",X"00",X"00",X"0F",X"3F",X"30",X"F0",
		X"00",X"00",X"03",X"FE",X"EE",X"F0",X"00",X"0E",X"F3",X"EE",X"EE",X"EF",X"00",X"00",X"03",X"EF",
		X"EE",X"57",X"F0",X"00",X"03",X"EF",X"EE",X"88",X"E0",X"0E",X"F3",X"EF",X"F7",X"88",X"70",X"00",
		X"03",X"EF",X"FF",X"57",X"F0",X"00",X"00",X"EF",X"F0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"00",X"0E",X"EF",X"EE",X"EE",X"00",X"00",X"EF",X"FE",X"EF",X"EE",X"E0",X"00",X"FF",X"0F",X"EF",
		X"3E",X"E0",X"00",X"0F",X"3F",X"EF",X"FE",X"E0",X"00",X"00",X"FE",X"EE",X"F0",X"EE",X"F0",X"00",
		X"FF",X"EE",X"EF",X"0E",X"E0",X"00",X"FF",X"0F",X"EE",X"0E",X"E0",X"00",X"EF",X"00",X"EE",X"0F",
		X"00",X"00",X"EE",X"00",X"EE",X"00",X"00",X"00",X"EE",X"E0",X"EE",X"00",X"00",X"00",X"EE",X"E0",
		X"EE",X"FE",X"00",X"00",X"FE",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",
		X"00",X"00",X"FE",X"00",X"00",X"0F",X"EE",X"EE",X"30",X"00",X"00",X"FE",X"EF",X"EE",X"E0",X"00",
		X"00",X"F2",X"EF",X"3E",X"F0",X"EE",X"00",X"0F",X"EF",X"FE",X"EE",X"EE",X"00",X"03",X"EE",X"FF",
		X"EF",X"F0",X"00",X"0F",X"3E",X"EF",X"3F",X"00",X"00",X"0E",X"F0",X"00",X"FE",X"00",X"00",X"0E",
		X"00",X"0F",X"EE",X"00",X"00",X"FE",X"00",X"0E",X"3E",X"F0",X"00",X"EF",X"E0",X"00",X"F3",X"E0",
		X"00",X"EE",X"E0",X"00",X"0F",X"E0",X"00",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"E0",X"EE",X"EE",X"00",X"00",X"00",X"0F",X"E0",X"FF",X"EE",X"00",
		X"00",X"00",X"0F",X"2E",X"EF",X"EE",X"00",X"00",X"00",X"00",X"FE",X"EF",X"EE",X"F0",X"00",X"00",
		X"00",X"0E",X"EF",X"EE",X"EE",X"00",X"00",X"00",X"0F",X"FE",X"FF",X"EF",X"E0",X"00",X"00",X"0F",
		X"F3",X"FF",X"FF",X"E0",X"00",X"00",X"0E",X"EF",X"00",X"0F",X"E0",X"00",X"EE",X"EE",X"F0",X"00",
		X"0E",X"FF",X"E0",X"FE",X"F0",X"00",X"00",X"0E",X"EE",X"F0",X"3E",X"F0",X"00",X"00",X"0E",X"EF",
		X"00",X"0E",X"E0",X"00",X"00",X"0F",X"E0",X"00",X"00",X"0F",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"E0",X"EE",X"EE",X"30",X"00",X"0F",X"FF",X"FE",X"EF",X"EE",X"E0",X"00",X"0F",X"F0",X"02",
		X"EF",X"3E",X"E0",X"00",X"0F",X"E0",X"0F",X"EF",X"FE",X"E0",X"E0",X"0E",X"F0",X"0E",X"EE",X"FF",
		X"EE",X"E0",X"00",X"00",X"00",X"EE",X"EF",X"8E",X"F0",X"00",X"00",X"EE",X"F8",X"EE",X"F0",X"00",
		X"00",X"00",X"E3",X"E3",X"EE",X"00",X"00",X"00",X"00",X"E3",X"E0",X"FE",X"00",X"00",X"00",X"00",
		X"0E",X"E0",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"0E",X"E0",X"EE",X"EE",X"00",X"00",X"00",X"0F",
		X"FE",X"EF",X"EE",X"E0",X"00",X"00",X"0F",X"02",X"EF",X"3E",X"E0",X"00",X"00",X"0F",X"F0",X"EF",
		X"FE",X"E0",X"EE",X"00",X"0F",X"E0",X"EE",X"FF",X"EE",X"EE",X"00",X"00",X"00",X"FE",X"EE",X"FF",
		X"0F",X"00",X"00",X"00",X"FF",X"8E",X"EE",X"00",X"00",X"00",X"00",X"0F",X"F0",X"0E",X"E0",X"00",
		X"00",X"00",X"0F",X"F0",X"EE",X"00",X"00",X"00",X"00",X"0F",X"EE",X"E0",X"00",X"00",X"00",X"00",
		X"0E",X"EE",X"00",X"00",X"00",X"00",X"00",X"03",X"E0",X"00",X"00",X"00",X"00",X"00",X"03",X"EF",
		X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"0E",X"E0",X"EE",X"FE",X"00",X"00",
		X"00",X"FE",X"FE",X"EF",X"EE",X"E0",X"00",X"00",X"FE",X"0F",X"FE",X"EE",X"F0",X"00",X"00",X"FF",
		X"00",X"FE",X"EF",X"00",X"00",X"00",X"0F",X"F3",X"FE",X"EE",X"EE",X"00",X"00",X"00",X"0E",X"FF",
		X"FF",X"EE",X"E0",X"00",X"00",X"0F",X"FE",X"EE",X"FF",X"F0",X"00",X"00",X"0F",X"F3",X"EE",X"EE",
		X"E0",X"00",X"00",X"00",X"EF",X"00",X"0E",X"E0",X"00",X"00",X"00",X"EE",X"00",X"0E",X"F0",X"00",
		X"00",X"FE",X"EF",X"00",X"0E",X"EE",X"00",X"00",X"F3",X"E0",X"00",X"0E",X"EF",X"00",X"00",X"F3",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"0F",X"E0",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"F0",X"EE",X"EE",X"30",X"00",X"00",X"00",X"FE",X"FF",X"FE",X"FE",
		X"EE",X"00",X"00",X"00",X"FF",X"00",X"FE",X"3E",X"EE",X"E0",X"00",X"00",X"FE",X"00",X"0E",X"F3",
		X"FE",X"EE",X"EE",X"F0",X"0E",X"F0",X"FE",X"EF",X"F0",X"00",X"EE",X"E0",X"0F",X"F0",X"EE",X"EE",
		X"F0",X"00",X"00",X"E0",X"0F",X"00",X"0E",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"EF",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"FE",X"EF",X"F0",X"00",X"00",X"00",X"00",X"0F",X"EE",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"FE",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"0E",X"00",X"F0",X"0E",X"00",X"00",X"F3",X"33",X"F0",X"00",X"00",X"33",X"FE",X"EE",X"50",
		X"EF",X"3F",X"EE",X"EE",X"80",X"03",X"3F",X"EF",X"E7",X"70",X"00",X"3F",X"EF",X"EE",X"50",X"EF",
		X"FF",X"EF",X"FE",X"00",X"00",X"3F",X"EF",X"00",X"00",X"00",X"3F",X"EF",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"EE",X"00",X"00",X"00",X"0E",X"FE",X"3E",X"E0",X"00",X"00",X"FF",X"EE",X"3E",X"E0",
		X"00",X"0F",X"EF",X"EF",X"FE",X"E0",X"00",X"EE",X"FF",X"FE",X"EE",X"00",X"0E",X"EF",X"0F",X"EE",
		X"FF",X"F0",X"0E",X"F0",X"0F",X"EE",X"FF",X"F0",X"00",X"E0",X"0F",X"EE",X"3E",X"E0",X"00",X"00",
		X"0E",X"FF",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"0E",X"F0",X"00",X"00",X"FE",X"E0",X"0E",X"E0",
		X"00",X"0F",X"EE",X"F0",X"0E",X"E0",X"00",X"0E",X"EF",X"00",X"FE",X"E0",X"00",X"00",X"00",X"0F",
		X"EE",X"F0",X"00",X"00",X"00",X"0E",X"EF",X"00",X"00",X"00",X"00",X"0F",X"EE",X"00",X"00",X"00",
		X"00",X"00",X"FE",X"3E",X"E0",X"00",X"00",X"0F",X"E3",X"FE",X"33",X"EE",X"00",X"EE",X"0E",X"FE",
		X"EE",X"F3",X"EE",X"00",X"EE",X"FE",X"3E",X"EF",X"FE",X"E0",X"00",X"FF",X"E0",X"3F",X"EE",X"FE",
		X"00",X"00",X"00",X"00",X"0E",X"EE",X"FE",X"F0",X"00",X"00",X"00",X"EE",X"EF",X"0F",X"E0",X"00",
		X"00",X"00",X"EE",X"F0",X"00",X"00",X"00",X"00",X"00",X"FE",X"EF",X"00",X"00",X"00",X"00",X"00",
		X"02",X"EE",X"F0",X"00",X"00",X"00",X"00",X"EF",X"FE",X"E0",X"00",X"00",X"00",X"0E",X"EF",X"EE",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"0F",X"EE",X"00",X"00",
		X"00",X"0F",X"FE",X"FF",X"E0",X"00",X"00",X"3F",X"EE",X"F3",X"EE",X"00",X"00",X"3E",X"EE",X"F0",
		X"FE",X"00",X"0E",X"3E",X"EE",X"F0",X"EE",X"00",X"0F",X"3E",X"EF",X"FF",X"EF",X"00",X"00",X"0E",
		X"EE",X"3E",X"E0",X"00",X"00",X"0F",X"EE",X"0F",X"E0",X"00",X"00",X"00",X"EE",X"F0",X"00",X"00",
		X"00",X"00",X"EE",X"FE",X"00",X"00",X"00",X"00",X"EE",X"FF",X"00",X"00",X"00",X"00",X"EE",X"F0",
		X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"EE",X"F0",X"00",X"00",X"00",X"0F",
		X"EE",X"F0",X"00",X"00",X"00",X"FE",X"EF",X"00",X"00",X"00",X"00",X"FE",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"EE",X"00",X"00",X"00",X"0F",X"FF",X"3E",X"E0",X"00",X"00",X"0F",X"EF",
		X"3E",X"E0",X"00",X"00",X"0E",X"EF",X"FE",X"F0",X"00",X"00",X"FE",X"FE",X"EE",X"30",X"00",X"FF",
		X"EF",X"EE",X"EF",X"F0",X"0F",X"EE",X"EF",X"EE",X"3F",X"E0",X"0E",X"EF",X"00",X"EE",X"0E",X"E0",
		X"00",X"EE",X"00",X"00",X"0E",X"E0",X"00",X"0E",X"E0",X"00",X"0E",X"F0",X"00",X"0E",X"EE",X"00",
		X"0E",X"E0",X"00",X"EE",X"F0",X"00",X"0E",X"E0",X"0F",X"EF",X"00",X"00",X"FE",X"E0",X"00",X"00",
		X"00",X"0F",X"EE",X"F0",X"00",X"00",X"00",X"0E",X"EF",X"00",X"00",X"00",X"00",X"FF",X"EE",X"00",
		X"00",X"00",X"00",X"0F",X"FE",X"3F",X"EE",X"00",X"00",X"00",X"3F",X"EE",X"F3",X"FE",X"E0",X"00",
		X"00",X"FE",X"EE",X"FE",X"EE",X"E0",X"0E",X"EF",X"3E",X"EE",X"EE",X"EF",X"00",X"0E",X"FF",X"3E",
		X"EE",X"3F",X"00",X"00",X"0E",X"00",X"EE",X"EE",X"F0",X"00",X"00",X"00",X"0E",X"EE",X"FE",X"E0",
		X"00",X"00",X"00",X"EE",X"E0",X"0E",X"E0",X"00",X"00",X"00",X"EE",X"00",X"0E",X"EF",X"EE",X"00",
		X"00",X"EF",X"00",X"0F",X"EE",X"FE",X"00",X"00",X"EE",X"00",X"00",X"0F",X"EE",X"00",X"0F",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"FE",X"EE",X"00",X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"EE",X"E0",X"00",X"00",X"00",X"FE",X"EE",X"EE",X"00",X"00",
		X"3F",X"EE",X"F0",X"FF",X"E0",X"00",X"3E",X"EE",X"00",X"0E",X"E0",X"00",X"3E",X"EF",X"30",X"EE",
		X"00",X"0F",X"3E",X"EF",X"3E",X"E0",X"00",X"0F",X"3E",X"EE",X"3E",X"EF",X"00",X"00",X"03",X"EE",
		X"00",X"FF",X"00",X"00",X"00",X"EE",X"F0",X"00",X"00",X"00",X"00",X"EE",X"3F",X"00",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"FE",X"E0",X"00",X"00",X"00",X"00",X"0E",X"EF",X"00",
		X"00",X"00",X"00",X"0F",X"EE",X"F0",X"00",X"00",X"00",X"0E",X"EE",X"00",X"00",X"00",X"00",X"0E",
		X"E0",X"00",X"00",X"00",X"00",X"03",X"FE",X"E0",X"00",X"00",X"00",X"03",X"FF",X"EE",X"EE",X"00",
		X"00",X"00",X"0F",X"EE",X"E3",X"FF",X"E0",X"00",X"EF",X"0E",X"EE",X"EF",X"00",X"FE",X"00",X"EE",
		X"3E",X"EE",X"EE",X"00",X"EE",X"00",X"00",X"0F",X"E3",X"EE",X"0F",X"E0",X"00",X"00",X"03",X"3E",
		X"EE",X"0E",X"E0",X"00",X"00",X"0F",X"EE",X"F0",X"0F",X"EE",X"00",X"00",X"0E",X"E3",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"EE",X"EE",X"EF",X"00",X"00",X"00",X"00",X"33",X"0F",X"EE",X"00",X"00",
		X"00",X"00",X"FE",X"0F",X"EE",X"00",X"00",X"00",X"0F",X"EE",X"0F",X"E0",X"00",X"00",X"00",X"0E",
		X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"E0",X"0F",X"00",X"E0",
		X"00",X"00",X"F0",X"3F",X"3F",X"00",X"00",X"00",X"FE",X"EE",X"F3",X"00",X"00",X"0F",X"EE",X"EE",
		X"E3",X"FE",X"00",X"F7",X"5E",X"EF",X"E3",X"00",X"00",X"E8",X"8E",X"EF",X"E3",X"00",X"00",X"78",
		X"87",X"FF",X"E3",X"FE",X"00",X"F7",X"5F",X"FF",X"E3",X"00",X"00",X"00",X"00",X"FF",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"EE",X"EF",X"EE",X"00",X"00",X"EE",X"EF",
		X"EE",X"FF",X"E0",X"00",X"EE",X"3F",X"EF",X"0F",X"F0",X"00",X"EE",X"FF",X"EF",X"3F",X"00",X"FE",
		X"E0",X"FE",X"EE",X"F0",X"00",X"EE",X"0F",X"EE",X"EF",X"F0",X"00",X"EE",X"0E",X"EF",X"0F",X"F0",
		X"00",X"0F",X"0E",X"E0",X"0F",X"E0",X"00",X"00",X"0E",X"E0",X"0E",X"E0",X"00",X"00",X"0E",X"E0",
		X"EE",X"E0",X"00",X"0E",X"FE",X"E0",X"EE",X"E0",X"00",X"0E",X"EE",X"E0",X"0E",X"F0",X"00",X"00",
		X"EE",X"E0",X"00",X"00",X"00",X"00",X"0E",X"F0",X"00",X"00",X"00",X"00",X"00",X"3E",X"EE",X"EF",
		X"00",X"00",X"00",X"EE",X"EF",X"EE",X"F0",X"0E",X"E0",X"FE",X"3F",X"E2",X"F0",X"0E",X"EE",X"EE",
		X"FF",X"EF",X"00",X"00",X"FF",X"EF",X"FE",X"E3",X"00",X"00",X"0F",X"3F",X"EE",X"3F",X"00",X"00",
		X"0E",X"F0",X"00",X"FE",X"00",X"00",X"0E",X"EF",X"00",X"0E",X"00",X"00",X"FE",X"3E",X"00",X"0E",
		X"F0",X"00",X"E3",X"F0",X"00",X"EF",X"E0",X"00",X"EF",X"00",X"00",X"EE",X"E0",X"00",X"00",X"00",
		X"00",X"0E",X"F0",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"0E",X"EE",X"E0",X"EE",
		X"00",X"00",X"00",X"0E",X"EF",X"F0",X"EF",X"00",X"00",X"00",X"0E",X"EF",X"EE",X"2F",X"00",X"00",
		X"00",X"FE",X"EF",X"EE",X"F0",X"00",X"00",X"0E",X"EE",X"EF",X"EE",X"00",X"00",X"00",X"EF",X"EF",
		X"FE",X"FF",X"00",X"00",X"00",X"EF",X"FF",X"F3",X"FF",X"00",X"00",X"00",X"EF",X"00",X"0F",X"EE",
		X"00",X"00",X"EF",X"FE",X"00",X"00",X"FE",X"EE",X"E0",X"FE",X"EE",X"00",X"00",X"00",X"FE",X"F0",
		X"0F",X"EE",X"00",X"00",X"00",X"FE",X"30",X"00",X"EF",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"00",X"00",X"EF",X"00",X"00",X"00",X"3E",X"EE",X"E0",X"EE",X"00",X"00",X"00",X"EE",X"EF",X"EE",
		X"FF",X"FF",X"00",X"00",X"EE",X"3F",X"E2",X"00",X"FF",X"00",X"E0",X"EE",X"FF",X"EF",X"00",X"EF",
		X"00",X"EE",X"EF",X"FE",X"EE",X"00",X"FE",X"00",X"FE",X"8F",X"EE",X"E0",X"00",X"00",X"00",X"00",
		X"FE",X"E8",X"FE",X"E0",X"00",X"00",X"00",X"0E",X"E3",X"E3",X"E0",X"00",X"00",X"00",X"0E",X"F0",
		X"E3",X"E0",X"00",X"00",X"00",X"0E",X"E0",X"EE",X"00",X"00",X"00",X"0E",X"FE",X"E0",X"00",X"00",
		X"00",X"00",X"0E",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"0E",X"EE",X"E0",X"EE",X"00",X"00",X"00",X"EE",X"EF",X"EE",X"FF",X"00",X"00",X"00",X"EE",X"3F",
		X"E2",X"0F",X"00",X"0E",X"E0",X"EE",X"FF",X"E0",X"FF",X"00",X"0E",X"EE",X"EF",X"FE",X"E0",X"EF",
		X"00",X"0F",X"0F",X"FE",X"EE",X"F0",X"00",X"00",X"00",X"0E",X"EE",X"8F",X"F0",X"00",X"00",X"00",
		X"EE",X"00",X"FF",X"00",X"00",X"00",X"00",X"0E",X"E0",X"FF",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"EF",X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"E3",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"E3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"0E",X"FE",X"E0",X"EE",X"00",X"00",X"00",X"EE",X"EF",X"EE",X"FE",X"F0",X"00",X"00",
		X"FE",X"EE",X"FF",X"0E",X"F0",X"00",X"00",X"0F",X"EE",X"F0",X"0F",X"F0",X"00",X"0E",X"EE",X"EE",
		X"F3",X"FF",X"00",X"00",X"EE",X"EF",X"FF",X"FE",X"00",X"00",X"00",X"FF",X"FE",X"EE",X"FF",X"00",
		X"00",X"00",X"EE",X"EE",X"E3",X"FF",X"00",X"00",X"00",X"EE",X"00",X"0F",X"E0",X"00",X"00",X"00",
		X"FE",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"EE",X"00",X"0F",X"EE",X"F0",X"00",X"0F",X"EE",X"00",
		X"00",X"E3",X"F0",X"00",X"00",X"00",X"00",X"00",X"E3",X"F0",X"00",X"00",X"00",X"00",X"00",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"3E",X"EE",X"E0",
		X"FE",X"00",X"00",X"00",X"0E",X"EE",X"FE",X"FF",X"FE",X"F0",X"00",X"00",X"EE",X"EE",X"3E",X"F0",
		X"0F",X"F0",X"FE",X"EE",X"EE",X"F3",X"FE",X"00",X"0E",X"F0",X"EE",X"E0",X"00",X"FF",X"EE",X"F0",
		X"FE",X"00",X"E0",X"00",X"00",X"FE",X"EE",X"E0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"EE",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"EF",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"EE",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"0E",X"E3",X"F0",X"00",X"00",X"00",X"00",X"00",X"0E",X"3F",
		X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"00",X"F0",X"0E",X"00",X"00",X"F3",X"33",X"F0",
		X"00",X"5E",X"EE",X"F3",X"30",X"00",X"8E",X"EE",X"EF",X"3F",X"E0",X"77",X"EF",X"EF",X"33",X"00",
		X"5E",X"EF",X"EF",X"30",X"00",X"0E",X"FF",X"EF",X"FF",X"E0",X"00",X"0F",X"EF",X"30",X"00",X"00",
		X"0F",X"EF",X"30",X"00",X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"00",
		X"88",X"88",X"88",X"00",X"00",X"08",X"00",X"00",X"08",X"00",X"00",X"08",X"00",X"00",X"08",X"00",
		X"88",X"88",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"08",
		X"88",X"80",X"08",X"00",X"00",X"08",X"00",X"00",X"08",X"00",X"00",X"08",X"88",X"88",X"80",X"08",
		X"88",X"88",X"80",X"08",X"88",X"88",X"80",X"08",X"88",X"88",X"80",X"08",X"00",X"00",X"08",X"00",
		X"00",X"08",X"00",X"00",X"08",X"00",X"00",X"08",X"88",X"80",X"00",X"00",X"80",X"00",X"00",X"00",
		X"80",X"00",X"00",X"80",X"00",X"00",X"88",X"88",X"00",X"00",X"08",X"00",X"00",X"08",X"00",X"00",
		X"08",X"00",X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"00",X"88",X"88",
		X"88",X"00",X"80",X"00",X"00",X"88",X"88",X"00",X"00",X"08",X"00",X"00",X"08",X"00",X"00",X"08",
		X"00",X"00",X"08",X"00",X"08",X"00",X"00",X"08",X"00",X"00",X"08",X"00",X"00",X"08",X"88",X"80",
		X"00",X"00",X"80",X"00",X"00",X"80",X"08",X"88",X"88",X"80",X"08",X"88",X"88",X"80",X"08",X"88",
		X"88",X"80",X"08",X"88",X"88",X"80",X"00",X"00",X"80",X"08",X"88",X"80",X"08",X"00",X"00",X"08",
		X"00",X"00",X"08",X"00",X"00",X"08",X"00",X"00",X"00",X"08",X"00",X"00",X"08",X"00",X"00",X"08",
		X"00",X"88",X"88",X"00",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"FE",X"FE",X"F0",X"00",
		X"00",X"00",X"0F",X"8F",X"EF",X"8F",X"00",X"00",X"00",X"FF",X"2F",X"EF",X"2F",X"F0",X"00",X"0F",
		X"F2",X"6F",X"EF",X"62",X"FF",X"00",X"02",X"F2",X"2F",X"EF",X"22",X"F2",X"00",X"F6",X"2F",X"3F",
		X"EF",X"3F",X"26",X"F0",X"2F",X"EE",X"8F",X"2F",X"8E",X"EF",X"20",X"22",X"FE",X"EF",X"2F",X"EE",
		X"F2",X"20",X"FE",X"EF",X"EF",X"2F",X"EF",X"EE",X"F0",X"2F",X"EE",X"FE",X"2E",X"FE",X"EF",X"20",
		X"62",X"FE",X"EF",X"6F",X"EE",X"F2",X"60",X"FE",X"EF",X"EE",X"6E",X"EF",X"EE",X"F0",X"2F",X"EE",
		X"FE",X"8E",X"FE",X"EF",X"20",X"FE",X"FE",X"EE",X"6E",X"EE",X"FE",X"F0",X"2F",X"DF",X"FE",X"8E",
		X"FF",X"DF",X"20",X"FE",X"FE",X"EE",X"6E",X"EE",X"FE",X"F0",X"2F",X"DF",X"FF",X"8F",X"FF",X"DF",
		X"20",X"FE",X"FE",X"EE",X"6E",X"EE",X"FE",X"F0",X"2F",X"DF",X"FF",X"8F",X"FF",X"DF",X"20",X"FE",
		X"FE",X"EE",X"6E",X"EE",X"FE",X"F0",X"2F",X"DF",X"FF",X"8F",X"FF",X"DF",X"20",X"FE",X"FE",X"EE",
		X"6E",X"EE",X"FE",X"F0",X"02",X"FD",X"FF",X"8F",X"FD",X"F2",X"00",X"00",X"FE",X"EE",X"6E",X"EE",
		X"F0",X"00",X"00",X"02",X"FF",X"8F",X"F2",X"00",X"00",X"00",X"00",X"0E",X"2E",X"00",X"00",X"00",
		X"10",X"11",X"10",X"11",X"10",X"11",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"11",
		X"10",X"11",X"10",X"11",X"10",X"00",X"00",X"00",X"A5",X"71",X"10",X"00",X"00",X"A5",X"77",X"71",
		X"A0",X"00",X"06",X"5A",X"00",X"75",X"00",X"0A",X"90",X"00",X"0A",X"70",X"00",X"00",X"00",X"00",
		X"05",X"00",X"00",X"11",X"75",X"A0",X"00",X"00",X"00",X"A1",X"77",X"75",X"A0",X"00",X"00",X"05",
		X"70",X"0A",X"56",X"00",X"00",X"00",X"7A",X"00",X"00",X"9A",X"00",X"00",X"05",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"0A",X"50",X"00",X"0A",X"60",X"00",X"00",X"06",X"7A",
		X"00",X"56",X"00",X"00",X"00",X"A5",X"77",X"71",X"A0",X"00",X"00",X"00",X"A5",X"71",X"10",X"00",
		X"0A",X"00",X"00",X"00",X"00",X"00",X"6A",X"00",X"00",X"5A",X"00",X"06",X"50",X"0A",X"76",X"00",
		X"00",X"A1",X"77",X"75",X"A0",X"00",X"00",X"11",X"75",X"A0",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
