library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity inferno_sound is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of inferno_sound is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"AD",X"0F",X"8E",X"00",X"7F",X"8D",X"02",X"20",X"FE",X"CE",X"20",X"00",X"6F",X"01",X"6F",X"03",
		X"86",X"FF",X"A7",X"02",X"C6",X"80",X"E7",X"00",X"86",X"37",X"A7",X"01",X"86",X"3C",X"A7",X"03",
		X"E7",X"00",X"0E",X"86",X"C6",X"97",X"64",X"39",X"7F",X"00",X"59",X"7F",X"00",X"5A",X"CE",X"EE",
		X"89",X"DF",X"6B",X"CE",X"EF",X"4B",X"DF",X"6D",X"BD",X"E7",X"F8",X"20",X"FE",X"BD",X"E7",X"80",
		X"BD",X"E7",X"B7",X"CE",X"00",X"00",X"DF",X"5E",X"7F",X"00",X"60",X"CE",X"00",X"20",X"DF",X"5C",
		X"7A",X"00",X"41",X"27",X"03",X"7E",X"E1",X"31",X"96",X"40",X"9B",X"59",X"9B",X"5A",X"97",X"41",
		X"DE",X"5E",X"A6",X"00",X"D6",X"45",X"27",X"10",X"D6",X"47",X"26",X"0C",X"16",X"54",X"27",X"03",
		X"54",X"26",X"02",X"C9",X"00",X"10",X"A7",X"00",X"B7",X"20",X"02",X"96",X"48",X"27",X"14",X"DE",
		X"5C",X"A6",X"00",X"16",X"C4",X"0F",X"44",X"44",X"44",X"44",X"DB",X"60",X"24",X"03",X"7C",X"00",
		X"5F",X"D7",X"60",X"9B",X"5F",X"4C",X"94",X"72",X"97",X"5F",X"27",X"03",X"7E",X"E1",X"31",X"DE",
		X"6D",X"A6",X"0E",X"27",X"0A",X"D6",X"65",X"7C",X"00",X"65",X"11",X"27",X"02",X"20",X"39",X"7F",
		X"00",X"65",X"A6",X"0F",X"2B",X"11",X"27",X"0A",X"D6",X"66",X"7C",X"00",X"66",X"11",X"27",X"02",
		X"20",X"26",X"7F",X"00",X"66",X"20",X"FE",X"84",X"7F",X"27",X"0A",X"D6",X"66",X"5C",X"11",X"27",
		X"04",X"D7",X"66",X"20",X"13",X"EE",X"10",X"DF",X"6D",X"BD",X"E7",X"F8",X"7F",X"00",X"66",X"7F",
		X"00",X"59",X"7F",X"00",X"5A",X"7E",X"E0",X"3D",X"96",X"54",X"27",X"05",X"7A",X"00",X"55",X"26",
		X"2C",X"DE",X"6B",X"A6",X"01",X"97",X"54",X"97",X"55",X"27",X"1A",X"A6",X"00",X"97",X"40",X"97",
		X"41",X"A6",X"02",X"97",X"42",X"97",X"43",X"08",X"08",X"08",X"DF",X"6B",X"7F",X"00",X"59",X"7F",
		X"00",X"5A",X"7E",X"E0",X"3D",X"A6",X"00",X"2C",X"FE",X"EE",X"03",X"DF",X"6B",X"D6",X"45",X"27",
		X"10",X"96",X"47",X"26",X"09",X"96",X"46",X"97",X"47",X"5A",X"D7",X"45",X"20",X"03",X"4A",X"97",
		X"47",X"96",X"48",X"27",X"4B",X"7A",X"00",X"49",X"26",X"46",X"97",X"49",X"D6",X"4D",X"27",X"1D",
		X"D6",X"4F",X"26",X"19",X"DE",X"5C",X"A6",X"00",X"16",X"54",X"27",X"0C",X"54",X"27",X"09",X"54",
		X"27",X"06",X"54",X"27",X"03",X"54",X"26",X"02",X"C9",X"00",X"10",X"A7",X"00",X"DE",X"5C",X"96",
		X"5D",X"4C",X"97",X"5D",X"81",X"40",X"26",X"18",X"80",X"20",X"97",X"5D",X"D6",X"4D",X"27",X"10",
		X"D6",X"4F",X"27",X"05",X"5A",X"D7",X"4F",X"20",X"07",X"D6",X"4E",X"D7",X"4F",X"7A",X"00",X"4D",
		X"96",X"58",X"85",X"01",X"27",X"2F",X"7A",X"00",X"51",X"26",X"2D",X"16",X"CE",X"00",X"59",X"C4",
		X"0C",X"27",X"15",X"C1",X"04",X"26",X"05",X"CE",X"00",X"44",X"20",X"0C",X"C1",X"08",X"26",X"05",
		X"CE",X"00",X"48",X"20",X"03",X"CE",X"00",X"4C",X"A6",X"00",X"94",X"57",X"4C",X"A7",X"00",X"D6",
		X"50",X"D7",X"51",X"20",X"03",X"7F",X"00",X"59",X"96",X"58",X"85",X"02",X"26",X"06",X"7F",X"00",
		X"5A",X"7E",X"E0",X"50",X"7A",X"00",X"53",X"26",X"44",X"D6",X"52",X"D7",X"53",X"4D",X"2B",X"08",
		X"CE",X"00",X"59",X"7F",X"00",X"5A",X"20",X"03",X"CE",X"00",X"5A",X"84",X"0C",X"27",X"15",X"81",
		X"04",X"26",X"05",X"CE",X"00",X"42",X"20",X"0C",X"81",X"08",X"26",X"05",X"CE",X"00",X"48",X"20",
		X"03",X"CE",X"00",X"4A",X"A6",X"00",X"81",X"01",X"22",X"03",X"7F",X"00",X"5B",X"91",X"56",X"23",
		X"03",X"7C",X"00",X"5B",X"4C",X"D6",X"5B",X"27",X"02",X"80",X"02",X"A7",X"00",X"7E",X"E0",X"50",
		X"96",X"4E",X"84",X"0F",X"27",X"1E",X"81",X"01",X"26",X"03",X"7E",X"E3",X"80",X"81",X"02",X"26",
		X"03",X"7E",X"E2",X"B8",X"81",X"03",X"26",X"03",X"7E",X"E3",X"2D",X"81",X"04",X"26",X"03",X"7E",
		X"E2",X"7B",X"20",X"FE",X"BD",X"E8",X"80",X"96",X"4A",X"B7",X"20",X"02",X"BD",X"E9",X"47",X"96",
		X"40",X"4A",X"26",X"FD",X"B6",X"20",X"02",X"16",X"54",X"54",X"54",X"10",X"7A",X"00",X"43",X"26",
		X"FA",X"9B",X"4B",X"D6",X"42",X"D7",X"43",X"B7",X"20",X"02",X"7A",X"00",X"47",X"26",X"07",X"7C",
		X"00",X"4B",X"96",X"46",X"97",X"47",X"7A",X"00",X"45",X"26",X"D1",X"7C",X"00",X"4A",X"96",X"44",
		X"97",X"45",X"BD",X"E8",X"D6",X"27",X"C0",X"2A",X"97",X"20",X"FE",X"96",X"4A",X"B7",X"20",X"02",
		X"BD",X"E9",X"47",X"96",X"40",X"4A",X"26",X"FD",X"B6",X"20",X"02",X"16",X"54",X"54",X"54",X"10",
		X"7A",X"00",X"43",X"26",X"FA",X"D6",X"42",X"D7",X"43",X"73",X"20",X"02",X"7A",X"00",X"45",X"26",
		X"0D",X"96",X"44",X"97",X"45",X"B6",X"20",X"02",X"BD",X"E8",X"68",X"B7",X"20",X"02",X"BD",X"E8",
		X"D6",X"27",X"CD",X"2B",X"FE",X"7E",X"E2",X"10",X"CE",X"00",X"00",X"7F",X"00",X"60",X"86",X"A5",
		X"C6",X"5A",X"97",X"61",X"D7",X"62",X"96",X"64",X"97",X"63",X"BD",X"E7",X"48",X"A7",X"00",X"A7",
		X"20",X"08",X"8C",X"00",X"20",X"26",X"F3",X"CE",X"00",X"00",X"C6",X"0C",X"86",X"80",X"A7",X"00",
		X"08",X"5A",X"26",X"FA",X"B7",X"20",X"02",X"BD",X"E9",X"47",X"CE",X"00",X"00",X"96",X"40",X"4A",
		X"26",X"FD",X"A6",X"01",X"AB",X"00",X"44",X"A7",X"00",X"B6",X"20",X"02",X"16",X"54",X"54",X"54",
		X"10",X"7A",X"00",X"43",X"26",X"FA",X"E6",X"00",X"54",X"1B",X"84",X"FC",X"D6",X"42",X"D7",X"43",
		X"B7",X"20",X"02",X"08",X"8C",X"00",X"3F",X"26",X"D4",X"A6",X"00",X"CE",X"00",X"00",X"AB",X"00",
		X"44",X"A7",X"3F",X"BD",X"E8",X"D6",X"27",X"BF",X"2B",X"FE",X"7E",X"E2",X"10",X"CE",X"00",X"00",
		X"7F",X"00",X"60",X"86",X"A5",X"C6",X"5A",X"97",X"61",X"D7",X"62",X"96",X"64",X"97",X"63",X"BD",
		X"E7",X"48",X"A7",X"00",X"08",X"8C",X"00",X"40",X"26",X"F5",X"7F",X"20",X"02",X"BD",X"E9",X"47",
		X"CE",X"00",X"00",X"96",X"40",X"4A",X"26",X"FD",X"B6",X"20",X"02",X"16",X"54",X"54",X"54",X"10",
		X"7A",X"00",X"43",X"26",X"FA",X"E6",X"00",X"54",X"1B",X"D6",X"42",X"D7",X"43",X"B7",X"20",X"02",
		X"08",X"8C",X"00",X"3F",X"26",X"DD",X"BD",X"E8",X"D6",X"27",X"D2",X"2B",X"FE",X"7E",X"E2",X"10",
		X"CE",X"00",X"00",X"86",X"FF",X"A7",X"00",X"08",X"8C",X"00",X"07",X"26",X"F8",X"7F",X"00",X"60",
		X"86",X"A5",X"C6",X"5A",X"97",X"61",X"D7",X"62",X"96",X"64",X"97",X"63",X"96",X"60",X"D6",X"61",
		X"53",X"C5",X"09",X"26",X"05",X"53",X"46",X"56",X"20",X"09",X"53",X"C5",X"09",X"26",X"02",X"27",
		X"F5",X"44",X"56",X"97",X"60",X"D7",X"61",X"A7",X"00",X"08",X"8C",X"00",X"3F",X"26",X"DD",X"BD",
		X"E9",X"47",X"CE",X"00",X"00",X"96",X"40",X"4A",X"26",X"FD",X"A6",X"01",X"D6",X"63",X"58",X"24",
		X"02",X"D8",X"64",X"D7",X"63",X"D4",X"4D",X"26",X"05",X"AB",X"00",X"44",X"A7",X"00",X"D6",X"63",
		X"58",X"24",X"02",X"D8",X"64",X"D7",X"63",X"D4",X"4C",X"27",X"03",X"40",X"A7",X"00",X"B6",X"20",
		X"02",X"16",X"54",X"54",X"54",X"10",X"7A",X"00",X"43",X"26",X"FA",X"E6",X"00",X"54",X"1B",X"84",
		X"FC",X"D6",X"42",X"D7",X"43",X"B7",X"20",X"02",X"08",X"8C",X"00",X"3F",X"26",X"B7",X"A6",X"00",
		X"CE",X"00",X"00",X"D6",X"63",X"58",X"24",X"02",X"D8",X"64",X"D7",X"63",X"D4",X"4D",X"26",X"05",
		X"AB",X"00",X"44",X"A7",X"3F",X"D6",X"63",X"58",X"24",X"02",X"D8",X"64",X"D7",X"63",X"D4",X"4C",
		X"27",X"01",X"40",X"B7",X"20",X"02",X"BD",X"E8",X"D6",X"27",X"84",X"2B",X"FE",X"7E",X"E2",X"10",
		X"BD",X"E9",X"83",X"CE",X"00",X"00",X"DF",X"6F",X"86",X"60",X"97",X"42",X"97",X"43",X"86",X"09",
		X"97",X"49",X"97",X"4A",X"7F",X"00",X"44",X"86",X"FF",X"97",X"47",X"96",X"40",X"4A",X"26",X"FD",
		X"DE",X"6F",X"E6",X"00",X"96",X"44",X"84",X"1F",X"BD",X"E7",X"64",X"EB",X"10",X"D4",X"47",X"F7",
		X"20",X"02",X"96",X"70",X"4C",X"97",X"70",X"81",X"40",X"26",X"E0",X"CE",X"00",X"00",X"DF",X"6F",
		X"96",X"48",X"27",X"1F",X"7A",X"00",X"4A",X"26",X"1A",X"D6",X"49",X"D7",X"4A",X"D6",X"40",X"C1",
		X"01",X"27",X"10",X"C1",X"25",X"27",X"0C",X"44",X"24",X"03",X"5A",X"20",X"04",X"44",X"24",X"03",
		X"5C",X"D7",X"40",X"7A",X"00",X"46",X"26",X"B3",X"7C",X"00",X"44",X"96",X"45",X"97",X"46",X"20",
		X"AA",X"16",X"58",X"1B",X"1B",X"1B",X"CE",X"FB",X"B2",X"BD",X"E7",X"64",X"A6",X"00",X"16",X"84",
		X"0F",X"97",X"0C",X"54",X"54",X"54",X"54",X"D7",X"0B",X"A6",X"01",X"16",X"54",X"54",X"54",X"54",
		X"D7",X"0D",X"84",X"0F",X"97",X"02",X"DF",X"04",X"CE",X"FA",X"EF",X"7A",X"00",X"02",X"2B",X"08",
		X"A6",X"00",X"4C",X"BD",X"E7",X"64",X"20",X"F3",X"DF",X"10",X"BD",X"E5",X"BC",X"DE",X"04",X"A6",
		X"02",X"97",X"12",X"9B",X"73",X"BD",X"E5",X"CE",X"7F",X"00",X"73",X"DE",X"04",X"A6",X"03",X"97",
		X"0E",X"A6",X"04",X"97",X"0F",X"A6",X"05",X"16",X"A6",X"06",X"CE",X"FC",X"06",X"BD",X"E7",X"64",
		X"17",X"DF",X"13",X"7F",X"00",X"1B",X"BD",X"E7",X"64",X"DF",X"15",X"39",X"96",X"0B",X"97",X"1A",
		X"DE",X"13",X"DF",X"06",X"DE",X"06",X"96",X"76",X"27",X"12",X"2B",X"10",X"DF",X"69",X"9B",X"6A",
		X"97",X"6A",X"5F",X"D9",X"69",X"D7",X"69",X"7F",X"00",X"76",X"DE",X"69",X"A6",X"00",X"9B",X"1B",
		X"97",X"19",X"9C",X"15",X"27",X"26",X"D6",X"0C",X"08",X"DF",X"06",X"CE",X"00",X"1C",X"96",X"19",
		X"4A",X"26",X"FD",X"A6",X"00",X"B7",X"20",X"02",X"08",X"9C",X"17",X"26",X"F1",X"5A",X"27",X"C4",
		X"08",X"09",X"08",X"09",X"08",X"09",X"08",X"09",X"01",X"01",X"20",X"DF",X"96",X"0D",X"8D",X"5E",
		X"7A",X"00",X"1A",X"26",X"AB",X"96",X"0E",X"27",X"42",X"7A",X"00",X"0F",X"27",X"3D",X"9B",X"1B",
		X"97",X"1B",X"DE",X"13",X"5F",X"96",X"1B",X"7D",X"00",X"0E",X"2B",X"06",X"AB",X"00",X"25",X"08",
		X"20",X"0B",X"AB",X"00",X"27",X"02",X"25",X"05",X"5D",X"27",X"08",X"20",X"0F",X"5D",X"26",X"03",
		X"DF",X"13",X"5C",X"08",X"9C",X"15",X"26",X"DD",X"5D",X"26",X"01",X"39",X"DF",X"15",X"96",X"0D",
		X"27",X"06",X"8D",X"08",X"96",X"12",X"8D",X"16",X"7E",X"E5",X"1C",X"39",X"CE",X"00",X"1C",X"DF",
		X"08",X"DE",X"10",X"E6",X"00",X"08",X"BD",X"E6",X"00",X"DE",X"08",X"DF",X"17",X"39",X"4D",X"27",
		X"2E",X"DE",X"10",X"DF",X"06",X"CE",X"00",X"1C",X"97",X"03",X"DF",X"08",X"DE",X"06",X"D6",X"03",
		X"D7",X"02",X"E6",X"01",X"54",X"54",X"54",X"54",X"08",X"DF",X"06",X"DE",X"08",X"A6",X"00",X"10",
		X"7A",X"00",X"02",X"26",X"FA",X"A7",X"00",X"08",X"9C",X"17",X"26",X"DE",X"7C",X"00",X"73",X"39",
		X"36",X"A6",X"00",X"DF",X"06",X"DE",X"08",X"A7",X"00",X"08",X"DF",X"08",X"DE",X"06",X"08",X"5A",
		X"26",X"EF",X"32",X"39",X"E6",X"1E",X"E6",X"23",X"01",X"01",X"01",X"FF",X"03",X"E8",X"CE",X"E6",
		X"18",X"20",X"07",X"4F",X"97",X"10",X"C6",X"03",X"20",X"10",X"A6",X"00",X"97",X"10",X"A6",X"01",
		X"97",X"11",X"A6",X"02",X"E6",X"03",X"EE",X"04",X"20",X"00",X"97",X"0F",X"D7",X"0A",X"DF",X"0D",
		X"7F",X"00",X"0C",X"86",X"AF",X"B7",X"20",X"02",X"97",X"00",X"97",X"01",X"DE",X"0D",X"B6",X"20",
		X"02",X"16",X"54",X"54",X"54",X"D8",X"01",X"54",X"76",X"00",X"00",X"76",X"00",X"01",X"D6",X"0A",
		X"7D",X"00",X"10",X"27",X"04",X"D4",X"00",X"DB",X"11",X"D7",X"0B",X"D6",X"0C",X"91",X"01",X"22",
		X"12",X"09",X"27",X"26",X"B7",X"20",X"02",X"DB",X"0C",X"99",X"0B",X"25",X"16",X"91",X"01",X"23",
		X"F0",X"20",X"10",X"09",X"27",X"14",X"B7",X"20",X"02",X"D0",X"0C",X"92",X"0B",X"25",X"04",X"91",
		X"01",X"22",X"F0",X"96",X"01",X"B7",X"20",X"02",X"20",X"B7",X"D6",X"0F",X"27",X"B3",X"96",X"0A",
		X"D6",X"0C",X"44",X"56",X"44",X"56",X"44",X"56",X"43",X"50",X"82",X"FF",X"DB",X"0C",X"99",X"0A",
		X"D7",X"0C",X"97",X"0A",X"26",X"96",X"C1",X"07",X"26",X"92",X"39",X"DE",X"6D",X"86",X"FF",X"B7",
		X"20",X"02",X"08",X"08",X"08",X"08",X"08",X"A6",X"03",X"97",X"03",X"A6",X"04",X"B7",X"20",X"02",
		X"A6",X"01",X"97",X"02",X"E6",X"00",X"2A",X"0F",X"C5",X"7F",X"27",X"FE",X"86",X"FF",X"4A",X"26",
		X"FD",X"5A",X"26",X"F8",X"08",X"20",X"E0",X"D7",X"01",X"A6",X"02",X"97",X"00",X"5A",X"26",X"FD",
		X"73",X"20",X"02",X"D6",X"01",X"4A",X"26",X"F5",X"96",X"00",X"DB",X"03",X"D7",X"01",X"D1",X"02",
		X"26",X"EB",X"20",X"BE",X"2A",X"1B",X"32",X"FF",X"FF",X"D8",X"2E",X"1D",X"22",X"FF",X"FF",X"23",
		X"49",X"0F",X"01",X"FF",X"80",X"2A",X"1B",X"32",X"FF",X"FF",X"D8",X"2E",X"1D",X"22",X"FF",X"FF",
		X"23",X"41",X"0F",X"01",X"FF",X"80",X"2D",X"0D",X"20",X"FF",X"FF",X"D8",X"30",X"19",X"22",X"FF",
		X"FF",X"19",X"47",X"0C",X"01",X"FF",X"80",X"49",X"31",X"12",X"FF",X"FF",X"D8",X"53",X"3A",X"15",
		X"FF",X"FF",X"38",X"61",X"10",X"01",X"FF",X"80",X"96",X"60",X"D6",X"61",X"53",X"C5",X"09",X"26",
		X"05",X"53",X"46",X"56",X"20",X"09",X"53",X"C5",X"09",X"26",X"02",X"27",X"F5",X"44",X"56",X"97",
		X"60",X"D7",X"61",X"39",X"DF",X"69",X"9B",X"6A",X"97",X"6A",X"96",X"69",X"89",X"00",X"97",X"69",
		X"DE",X"69",X"39",X"DF",X"69",X"DB",X"6A",X"D7",X"6A",X"99",X"69",X"97",X"69",X"DE",X"69",X"39",
		X"CE",X"00",X"00",X"DF",X"5E",X"DE",X"6F",X"DF",X"69",X"DE",X"69",X"A6",X"00",X"08",X"DF",X"69",
		X"D6",X"42",X"27",X"17",X"D7",X"67",X"16",X"54",X"27",X"09",X"54",X"27",X"06",X"54",X"27",X"03",
		X"54",X"26",X"02",X"C9",X"00",X"10",X"7A",X"00",X"67",X"26",X"EB",X"DE",X"5E",X"A7",X"00",X"7C",
		X"00",X"5F",X"9C",X"71",X"26",X"D3",X"39",X"CE",X"00",X"20",X"DF",X"5C",X"CE",X"ED",X"2A",X"DF",
		X"69",X"DE",X"69",X"A6",X"00",X"08",X"8C",X"ED",X"4A",X"26",X"03",X"CE",X"ED",X"2A",X"DF",X"69",
		X"D6",X"4A",X"27",X"17",X"D7",X"4B",X"16",X"54",X"27",X"09",X"54",X"27",X"06",X"54",X"27",X"03",
		X"54",X"26",X"02",X"C9",X"00",X"10",X"7A",X"00",X"4B",X"26",X"EB",X"DE",X"5C",X"A7",X"00",X"7C",
		X"00",X"5D",X"8C",X"00",X"3F",X"26",X"CA",X"39",X"36",X"DE",X"6D",X"A6",X"00",X"97",X"40",X"97",
		X"41",X"A6",X"01",X"97",X"42",X"97",X"43",X"A6",X"02",X"97",X"44",X"97",X"45",X"A6",X"03",X"97",
		X"46",X"97",X"47",X"A6",X"04",X"97",X"48",X"97",X"49",X"A6",X"05",X"97",X"4A",X"97",X"4B",X"A6",
		X"06",X"97",X"4C",X"97",X"4D",X"A6",X"07",X"97",X"4E",X"97",X"4F",X"A6",X"08",X"97",X"50",X"97",
		X"51",X"A6",X"09",X"97",X"52",X"97",X"53",X"A6",X"0A",X"97",X"54",X"97",X"55",X"A6",X"0B",X"97",
		X"56",X"A6",X"0C",X"97",X"57",X"A6",X"0D",X"97",X"58",X"85",X"10",X"26",X"19",X"DE",X"6B",X"A6",
		X"00",X"97",X"40",X"97",X"41",X"A6",X"01",X"97",X"54",X"97",X"55",X"A6",X"02",X"97",X"42",X"97",
		X"43",X"08",X"08",X"08",X"DF",X"6B",X"32",X"39",X"91",X"50",X"22",X"03",X"7F",X"00",X"52",X"91",
		X"51",X"23",X"03",X"7C",X"00",X"52",X"4C",X"D6",X"52",X"27",X"02",X"80",X"02",X"97",X"53",X"39",
		X"DE",X"6B",X"A6",X"00",X"97",X"40",X"97",X"41",X"A6",X"01",X"97",X"48",X"97",X"49",X"DE",X"6D",
		X"A6",X"01",X"97",X"42",X"97",X"43",X"A6",X"02",X"97",X"44",X"97",X"45",X"A6",X"03",X"97",X"46",
		X"97",X"47",X"A6",X"05",X"97",X"4A",X"A6",X"06",X"97",X"4B",X"A6",X"07",X"97",X"4C",X"A6",X"08",
		X"97",X"4D",X"A6",X"0A",X"97",X"4F",X"A6",X"09",X"97",X"4E",X"85",X"20",X"27",X"07",X"BD",X"E7",
		X"48",X"97",X"4A",X"96",X"4E",X"85",X"10",X"27",X"0C",X"A6",X"00",X"97",X"40",X"97",X"41",X"A6",
		X"04",X"97",X"48",X"97",X"49",X"39",X"DE",X"6D",X"A6",X"0B",X"27",X"0A",X"D6",X"65",X"5C",X"11",
		X"27",X"04",X"D7",X"65",X"20",X"32",X"7F",X"00",X"65",X"A6",X"0C",X"2B",X"11",X"27",X"0A",X"D6",
		X"66",X"7C",X"00",X"66",X"11",X"27",X"02",X"20",X"1F",X"7F",X"00",X"66",X"20",X"46",X"84",X"7F",
		X"27",X"0A",X"D6",X"66",X"5C",X"11",X"27",X"04",X"D7",X"66",X"20",X"0C",X"EE",X"0D",X"DF",X"6D",
		X"BD",X"E8",X"80",X"7F",X"00",X"66",X"20",X"29",X"96",X"48",X"27",X"05",X"7A",X"00",X"49",X"26",
		X"1E",X"DE",X"6B",X"A6",X"01",X"97",X"48",X"97",X"49",X"27",X"0C",X"A6",X"00",X"97",X"40",X"08",
		X"08",X"DF",X"6B",X"20",X"0C",X"20",X"0D",X"A6",X"00",X"2C",X"FE",X"EE",X"02",X"DF",X"6B",X"4F",
		X"39",X"86",X"01",X"39",X"86",X"FF",X"39",X"96",X"4F",X"44",X"24",X"06",X"7C",X"00",X"40",X"7C",
		X"00",X"41",X"44",X"24",X"06",X"7C",X"00",X"42",X"7C",X"00",X"43",X"44",X"24",X"06",X"7C",X"00",
		X"44",X"7C",X"00",X"45",X"44",X"24",X"06",X"7C",X"00",X"46",X"7C",X"00",X"47",X"44",X"24",X"06",
		X"7C",X"00",X"48",X"7C",X"00",X"49",X"44",X"24",X"03",X"7C",X"00",X"4C",X"44",X"24",X"03",X"7C",
		X"00",X"4D",X"39",X"CE",X"00",X"00",X"7F",X"00",X"60",X"86",X"A5",X"C6",X"5A",X"97",X"61",X"D7",
		X"62",X"96",X"64",X"97",X"63",X"96",X"60",X"D6",X"61",X"53",X"C5",X"09",X"26",X"05",X"53",X"46",
		X"56",X"20",X"09",X"53",X"C5",X"09",X"26",X"02",X"27",X"F5",X"44",X"56",X"97",X"60",X"D7",X"61",
		X"A7",X"00",X"08",X"8C",X"00",X"3F",X"26",X"DD",X"39",X"8E",X"00",X"7F",X"B6",X"20",X"00",X"0E",
		X"81",X"6F",X"26",X"07",X"97",X"02",X"BD",X"E0",X"09",X"96",X"02",X"81",X"AF",X"22",X"02",X"8D",
		X"28",X"86",X"3C",X"B7",X"20",X"03",X"86",X"37",X"B7",X"20",X"01",X"20",X"FE",X"0F",X"8E",X"00",
		X"7F",X"4F",X"CE",X"FF",X"FF",X"5F",X"E9",X"00",X"09",X"8C",X"E0",X"00",X"26",X"F8",X"E1",X"00",
		X"26",X"FE",X"86",X"01",X"8D",X"03",X"20",X"E5",X"39",X"C6",X"3C",X"F7",X"20",X"01",X"C6",X"3F",
		X"F7",X"20",X"01",X"4D",X"27",X"F2",X"D6",X"76",X"CA",X"80",X"D7",X"76",X"D6",X"75",X"81",X"A0",
		X"26",X"0B",X"7F",X"00",X"74",X"7F",X"00",X"73",X"7F",X"00",X"76",X"20",X"55",X"81",X"A4",X"26",
		X"0E",X"D6",X"74",X"CB",X"05",X"D7",X"73",X"D6",X"76",X"C4",X"7F",X"D7",X"76",X"20",X"43",X"C1",
		X"A0",X"26",X"1B",X"97",X"75",X"D6",X"73",X"D7",X"74",X"96",X"07",X"90",X"14",X"D6",X"06",X"D0",
		X"13",X"56",X"1B",X"8A",X"80",X"97",X"76",X"96",X"75",X"7F",X"00",X"73",X"20",X"26",X"C1",X"A4",
		X"26",X"1D",X"97",X"75",X"D6",X"74",X"DB",X"73",X"D7",X"74",X"96",X"07",X"90",X"14",X"D6",X"06",
		X"D0",X"13",X"56",X"1B",X"8A",X"80",X"97",X"76",X"96",X"75",X"7F",X"00",X"73",X"20",X"05",X"7F",
		X"00",X"73",X"97",X"75",X"CE",X"EB",X"AC",X"4A",X"16",X"4F",X"58",X"89",X"00",X"BD",X"E7",X"73",
		X"A6",X"00",X"E6",X"01",X"48",X"CE",X"EB",X"96",X"BD",X"E7",X"64",X"EE",X"00",X"17",X"6E",X"00",
		X"BD",X"E4",X"B1",X"7E",X"E5",X"1C",X"CE",X"E6",X"14",X"48",X"BD",X"E7",X"64",X"EE",X"00",X"6E",
		X"00",X"CE",X"EA",X"DA",X"48",X"1B",X"BD",X"E7",X"64",X"A6",X"00",X"97",X"40",X"A6",X"01",X"97",
		X"45",X"97",X"46",X"A6",X"02",X"97",X"48",X"7E",X"E4",X"40",X"CE",X"EA",X"D2",X"DF",X"69",X"48",
		X"9B",X"6A",X"24",X"03",X"7C",X"00",X"69",X"97",X"6A",X"DE",X"69",X"EE",X"00",X"DF",X"6D",X"7E",
		X"E6",X"BB",X"E6",X"FF",X"E7",X"10",X"E7",X"21",X"E7",X"32",X"20",X"04",X"00",X"19",X"08",X"01",
		X"13",X"09",X"01",X"05",X"05",X"02",X"CE",X"F3",X"BB",X"20",X"0D",X"CE",X"F2",X"5B",X"20",X"08",
		X"CE",X"F2",X"7B",X"20",X"03",X"CE",X"F2",X"9B",X"BD",X"E7",X"48",X"C4",X"03",X"20",X"06",X"7E",
		X"E9",X"D1",X"CE",X"F2",X"BB",X"4F",X"58",X"89",X"00",X"48",X"58",X"89",X"00",X"48",X"58",X"89",
		X"00",X"BD",X"E7",X"73",X"8C",X"F3",X"EB",X"27",X"E6",X"A6",X"00",X"97",X"6B",X"A6",X"01",X"97",
		X"6C",X"A6",X"02",X"97",X"6D",X"A6",X"03",X"97",X"6E",X"A6",X"04",X"97",X"6F",X"A6",X"05",X"97",
		X"70",X"A6",X"06",X"97",X"71",X"A6",X"07",X"97",X"72",X"DE",X"6B",X"BD",X"E7",X"F8",X"7F",X"00",
		X"66",X"7F",X"00",X"65",X"7F",X"00",X"59",X"7F",X"00",X"5A",X"7E",X"E0",X"3D",X"BD",X"E7",X"48",
		X"84",X"03",X"48",X"CE",X"EB",X"5D",X"BD",X"E7",X"64",X"EE",X"00",X"20",X"1B",X"FA",X"DF",X"FA",
		X"E3",X"FA",X"E7",X"FA",X"EB",X"4F",X"58",X"89",X"00",X"48",X"58",X"89",X"00",X"CE",X"F9",X"B7",
		X"BD",X"E7",X"73",X"8C",X"FA",X"EF",X"27",X"87",X"A6",X"00",X"97",X"6B",X"A6",X"01",X"97",X"6C",
		X"A6",X"02",X"97",X"6D",X"A6",X"03",X"97",X"6E",X"A6",X"04",X"BD",X"E8",X"80",X"7F",X"00",X"66",
		X"7F",X"00",X"65",X"7E",X"E2",X"10",X"EA",X"90",X"EA",X"96",X"EB",X"02",X"EB",X"65",X"EA",X"A1",
		X"EA",X"EB",X"EA",X"F0",X"EA",X"F5",X"EB",X"4D",X"EA",X"E6",X"EA",X"BA",X"00",X"00",X"00",X"01",
		X"00",X"02",X"00",X"03",X"00",X"04",X"01",X"00",X"04",X"00",X"05",X"00",X"06",X"00",X"07",X"00",
		X"02",X"00",X"02",X"24",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"00",X"00",X"00",X"00",X"02",X"04",
		X"00",X"00",X"00",X"00",X"02",X"05",X"02",X"06",X"02",X"07",X"02",X"08",X"02",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"0A",X"02",X"0B",X"00",X"00",X"02",X"0C",X"02",X"0D",X"02",X"0E",
		X"00",X"00",X"00",X"00",X"02",X"0E",X"02",X"0F",X"02",X"10",X"02",X"11",X"02",X"12",X"02",X"11",
		X"00",X"00",X"02",X"14",X"00",X"00",X"02",X"15",X"02",X"16",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"17",X"02",X"18",X"02",X"19",X"02",X"15",X"02",X"16",X"03",X"00",X"03",X"01",X"03",X"02",
		X"03",X"03",X"03",X"04",X"03",X"05",X"03",X"06",X"03",X"07",X"03",X"08",X"03",X"09",X"03",X"0A",
		X"03",X"0B",X"03",X"0C",X"03",X"0D",X"03",X"0E",X"03",X"0F",X"03",X"10",X"03",X"11",X"03",X"12",
		X"03",X"13",X"03",X"14",X"03",X"15",X"03",X"16",X"03",X"17",X"03",X"18",X"03",X"19",X"03",X"1A",
		X"03",X"1B",X"03",X"1C",X"03",X"1D",X"03",X"1E",X"03",X"1F",X"03",X"20",X"03",X"21",X"03",X"22",
		X"03",X"23",X"03",X"24",X"03",X"26",X"03",X"27",X"03",X"28",X"03",X"2A",X"03",X"2B",X"03",X"2F",
		X"03",X"30",X"03",X"31",X"03",X"32",X"03",X"33",X"03",X"34",X"03",X"35",X"03",X"36",X"03",X"37",
		X"03",X"38",X"03",X"39",X"04",X"01",X"04",X"02",X"00",X"05",X"00",X"06",X"01",X"01",X"02",X"17",
		X"03",X"3A",X"03",X"3B",X"03",X"3C",X"03",X"3D",X"03",X"3E",X"03",X"3F",X"03",X"40",X"03",X"41",
		X"03",X"42",X"03",X"43",X"03",X"44",X"03",X"45",X"03",X"46",X"03",X"47",X"02",X"18",X"02",X"1F",
		X"02",X"20",X"02",X"1B",X"02",X"22",X"02",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"48",X"03",X"49",X"08",X"00",X"03",X"4A",
		X"03",X"4B",X"03",X"4C",X"03",X"4D",X"02",X"24",X"00",X"00",X"00",X"07",X"00",X"08",X"00",X"09",
		X"00",X"0A",X"00",X"0B",X"09",X"00",X"02",X"20",X"02",X"21",X"02",X"22",X"02",X"23",X"0A",X"00",
		X"0A",X"01",X"0A",X"02",X"0A",X"03",X"04",X"03",X"02",X"25",X"99",X"B1",X"C8",X"DB",X"EB",X"F7",
		X"FE",X"FF",X"FE",X"F7",X"EB",X"DB",X"C8",X"B1",X"99",X"81",X"68",X"50",X"39",X"26",X"16",X"0A",
		X"03",X"01",X"03",X"0A",X"16",X"26",X"39",X"50",X"68",X"81",X"99",X"B1",X"C8",X"DB",X"EB",X"F7",
		X"FE",X"FF",X"FE",X"F7",X"EB",X"DB",X"C8",X"B1",X"99",X"81",X"68",X"50",X"39",X"26",X"16",X"0A",
		X"03",X"01",X"03",X"0A",X"16",X"26",X"39",X"50",X"68",X"81",X"B1",X"A8",X"B5",X"E7",X"F2",X"EC",
		X"FD",X"FE",X"FF",X"FE",X"E2",X"CD",X"D8",X"BA",X"81",X"81",X"80",X"47",X"29",X"34",X"1F",X"03",
		X"02",X"03",X"04",X"15",X"0F",X"1A",X"4C",X"59",X"50",X"81",X"DA",X"FA",X"FC",X"F4",X"ED",X"F6",
		X"FF",X"FC",X"FB",X"FF",X"E0",X"AA",X"9A",X"B8",X"DF",X"F1",X"EE",X"E0",X"DB",X"F4",X"FD",X"BF",
		X"76",X"5E",X"6E",X"84",X"7D",X"56",X"2D",X"20",X"3B",X"81",X"C6",X"E1",X"D4",X"AB",X"84",X"7D",
		X"93",X"A3",X"8B",X"42",X"04",X"0D",X"26",X"21",X"13",X"10",X"22",X"49",X"67",X"57",X"21",X"01",
		X"06",X"05",X"01",X"0B",X"14",X"0D",X"05",X"07",X"27",X"81",X"FB",X"FD",X"C5",X"A5",X"DF",X"FD",
		X"FC",X"FB",X"FF",X"EE",X"F5",X"FB",X"CA",X"3F",X"1E",X"81",X"E3",X"C2",X"37",X"06",X"0C",X"13",
		X"02",X"06",X"05",X"04",X"22",X"5C",X"3C",X"04",X"06",X"81",X"B9",X"B0",X"A4",X"94",X"80",X"6C",
		X"59",X"49",X"40",X"38",X"38",X"3A",X"3E",X"40",X"41",X"43",X"45",X"4B",X"53",X"5D",X"6B",X"7B",
		X"8F",X"9F",X"AF",X"B8",X"C5",X"CF",X"DB",X"E2",X"E2",X"DA",X"D0",X"C6",X"00",X"00",X"FF",X"00",
		X"ED",X"EE",X"04",X"04",X"04",X"1E",X"00",X"00",X"60",X"04",X"60",X"08",X"60",X"18",X"00",X"00",
		X"01",X"20",X"02",X"20",X"03",X"1D",X"02",X"20",X"04",X"10",X"03",X"20",X"05",X"0A",X"01",X"40",
		X"00",X"00",X"C0",X"07",X"C0",X"20",X"80",X"20",X"70",X"40",X"50",X"60",X"40",X"80",X"30",X"A0",
		X"20",X"C0",X"10",X"D0",X"FF",X"00",X"EE",X"12",X"09",X"C0",X"0A",X"BC",X"09",X"C0",X"0A",X"BC",
		X"09",X"C0",X"00",X"00",X"01",X"10",X"02",X"03",X"01",X"72",X"01",X"00",X"50",X"60",X"40",X"80",
		X"20",X"C0",X"10",X"D0",X"FF",X"00",X"EE",X"3C",X"01",X"2E",X"02",X"37",X"03",X"A1",X"04",X"EF",
		X"07",X"E6",X"00",X"00",X"03",X"2E",X"01",X"37",X"03",X"8B",X"04",X"8C",X"0B",X"72",X"10",X"FF",
		X"00",X"00",X"01",X"13",X"04",X"09",X"05",X"09",X"05",X"07",X"04",X"09",X"09",X"0F",X"09",X"0F",
		X"09",X"0F",X"01",X"10",X"04",X"09",X"03",X"07",X"05",X"09",X"04",X"09",X"09",X"0F",X"09",X"0F",
		X"09",X"0F",X"09",X"0F",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"EE",X"89",X"02",X"20",
		X"00",X"04",X"20",X"03",X"07",X"20",X"01",X"06",X"20",X"09",X"05",X"20",X"05",X"03",X"20",X"01",
		X"05",X"20",X"09",X"04",X"02",X"03",X"01",X"06",X"09",X"04",X"02",X"05",X"01",X"06",X"00",X"04",
		X"02",X"00",X"01",X"06",X"04",X"05",X"20",X"05",X"01",X"20",X"02",X"04",X"20",X"02",X"01",X"20",
		X"01",X"02",X"20",X"09",X"04",X"20",X"09",X"07",X"20",X"03",X"05",X"20",X"04",X"09",X"20",X"02",
		X"08",X"24",X"00",X"0A",X"09",X"01",X"0B",X"F0",X"00",X"00",X"00",X"00",X"06",X"07",X"00",X"07",
		X"07",X"00",X"08",X"05",X"00",X"00",X"00",X"00",X"00",X"07",X"02",X"00",X"06",X"04",X"00",X"05",
		X"18",X"00",X"00",X"00",X"00",X"08",X"02",X"00",X"07",X"04",X"00",X"06",X"0B",X"00",X"00",X"00",
		X"00",X"06",X"0B",X"00",X"07",X"04",X"00",X"04",X"10",X"00",X"00",X"00",X"00",X"01",X"03",X"00",
		X"04",X"10",X"00",X"00",X"00",X"00",X"05",X"07",X"02",X"03",X"1C",X"15",X"00",X"00",X"00",X"07",
		X"18",X"00",X"00",X"00",X"00",X"04",X"2C",X"00",X"00",X"00",X"00",X"01",X"28",X"00",X"02",X"27",
		X"00",X"03",X"26",X"00",X"06",X"1C",X"00",X"09",X"40",X"00",X"00",X"00",X"00",X"04",X"20",X"00",
		X"05",X"20",X"00",X"04",X"20",X"00",X"03",X"20",X"00",X"EF",X"3D",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"01",X"FF",X"20",X"0F",X"10",X"7F",X"FF",X"EF",X"4B",X"00",X"08",X"00",
		X"00",X"1F",X"05",X"00",X"00",X"15",X"05",X"FF",X"20",X"0F",X"11",X"FF",X"FF",X"EF",X"5D",X"00",
		X"08",X"00",X"00",X"1A",X"05",X"00",X"00",X"15",X"05",X"FF",X"20",X"0F",X"11",X"FF",X"FF",X"EF",
		X"6F",X"00",X"08",X"00",X"00",X"2B",X"05",X"00",X"00",X"15",X"05",X"FF",X"20",X"0F",X"11",X"FF",
		X"FF",X"EF",X"81",X"01",X"00",X"05",X"19",X"F4",X"00",X"00",X"00",X"0B",X"01",X"1B",X"10",X"0F",
		X"12",X"19",X"00",X"00",X"00",X"05",X"19",X"F4",X"00",X"00",X"00",X"0B",X"01",X"34",X"10",X"0F",
		X"12",X"31",X"00",X"FD",X"04",X"00",X"00",X"0D",X"13",X"00",X"00",X"0D",X"FA",X"FF",X"20",X"0F",
		X"91",X"FF",X"FF",X"EF",X"B3",X"FE",X"04",X"50",X"01",X"14",X"00",X"00",X"00",X"0D",X"FA",X"6E",
		X"20",X"0F",X"91",X"FF",X"00",X"05",X"00",X"51",X"19",X"DD",X"00",X"F3",X"00",X"FF",X"01",X"00",
		X"10",X"0F",X"00",X"FF",X"00",X"02",X"00",X"00",X"00",X"F4",X"00",X"0C",X"06",X"50",X"FC",X"00",
		X"21",X"0F",X"91",X"12",X"00",X"0A",X"01",X"00",X"00",X"01",X"07",X"00",X"00",X"03",X"09",X"FF",
		X"0F",X"0F",X"12",X"FF",X"FF",X"EF",X"F5",X"F9",X"00",X"1C",X"12",X"FF",X"00",X"E6",X"09",X"0D",
		X"1C",X"55",X"16",X"15",X"F3",X"09",X"80",X"F0",X"19",X"0A",X"10",X"00",X"00",X"01",X"07",X"00",
		X"00",X"03",X"09",X"FF",X"0F",X"0F",X"12",X"FF",X"7F",X"05",X"01",X"00",X"00",X"01",X"02",X"00",
		X"00",X"09",X"1F",X"FF",X"0F",X"0F",X"12",X"7F",X"75",X"0A",X"01",X"00",X"00",X"01",X"0F",X"00",
		X"00",X"09",X"1F",X"03",X"0F",X"0F",X"12",X"01",X"75",X"00",X"00",X"50",X"01",X"17",X"06",X"00",
		X"00",X"00",X"FF",X"09",X"20",X"0F",X"91",X"03",X"10",X"02",X"00",X"00",X"00",X"01",X"09",X"00",
		X"00",X"08",X"00",X"00",X"20",X"0F",X"00",X"10",X"81",X"02",X"00",X"00",X"00",X"01",X"05",X"00",
		X"00",X"08",X"00",X"00",X"20",X"0F",X"00",X"10",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"02",X"01",X"00",X"0F",X"0F",X"11",X"FF",X"00",X"01",X"00",X"80",X"09",X"00",X"00",X"00",
		X"00",X"02",X"01",X"00",X"0F",X"0F",X"10",X"FF",X"FF",X"F0",X"89",X"08",X"10",X"00",X"00",X"01",
		X"07",X"00",X"00",X"09",X"1F",X"FF",X"0F",X"00",X"12",X"FF",X"7F",X"12",X"0C",X"00",X"00",X"02",
		X"04",X"00",X"00",X"09",X"1F",X"FF",X"0F",X"0F",X"14",X"FF",X"7F",X"F9",X"00",X"1C",X"12",X"FF",
		X"00",X"E6",X"09",X"0D",X"1C",X"55",X"16",X"15",X"F3",X"1C",X"00",X"F9",X"00",X"1C",X"12",X"FF",
		X"00",X"E6",X"09",X"0D",X"1C",X"55",X"16",X"15",X"F3",X"1A",X"00",X"01",X"00",X"1C",X"12",X"F2",
		X"00",X"E8",X"08",X"0D",X"1C",X"55",X"16",X"15",X"13",X"32",X"00",X"01",X"00",X"1C",X"12",X"F2",
		X"00",X"E8",X"08",X"0D",X"1C",X"55",X"16",X"15",X"11",X"38",X"00",X"00",X"00",X"1C",X"12",X"F2",
		X"00",X"E8",X"08",X"0D",X"1C",X"55",X"16",X"15",X"11",X"38",X"00",X"02",X"00",X"00",X"00",X"02",
		X"02",X"80",X"03",X"0D",X"20",X"4A",X"13",X"13",X"1B",X"A9",X"00",X"01",X"00",X"1C",X"12",X"F2",
		X"00",X"E8",X"08",X"0D",X"1C",X"55",X"16",X"15",X"1C",X"4F",X"00",X"01",X"00",X"1C",X"12",X"F2",
		X"00",X"E8",X"08",X"0D",X"1C",X"55",X"16",X"15",X"1A",X"63",X"00",X"01",X"00",X"1C",X"12",X"F2",
		X"00",X"E8",X"08",X"0D",X"1C",X"55",X"16",X"15",X"18",X"73",X"00",X"01",X"00",X"1C",X"12",X"F2",
		X"00",X"E8",X"08",X"0D",X"1C",X"55",X"16",X"15",X"17",X"4D",X"00",X"00",X"02",X"1C",X"12",X"CD",
		X"13",X"DF",X"F4",X"35",X"0F",X"48",X"11",X"23",X"F1",X"9B",X"00",X"01",X"00",X"00",X"00",X"FF",
		X"08",X"26",X"13",X"0D",X"21",X"4A",X"14",X"15",X"13",X"2E",X"00",X"01",X"00",X"00",X"00",X"FF",
		X"06",X"26",X"13",X"0D",X"21",X"4A",X"14",X"0C",X"F1",X"3A",X"00",X"00",X"07",X"00",X"00",X"07",
		X"16",X"DF",X"F4",X"35",X"0F",X"48",X"11",X"23",X"F1",X"30",X"00",X"00",X"07",X"00",X"00",X"06",
		X"16",X"DF",X"F4",X"35",X"0F",X"48",X"11",X"23",X"F1",X"2E",X"00",X"01",X"07",X"00",X"00",X"3E",
		X"05",X"BA",X"10",X"34",X"0D",X"45",X"0F",X"19",X"F1",X"21",X"00",X"01",X"07",X"00",X"00",X"3C",
		X"0E",X"BA",X"F3",X"34",X"0D",X"45",X"0F",X"19",X"F1",X"1A",X"00",X"03",X"00",X"00",X"00",X"01",
		X"0E",X"00",X"00",X"04",X"1F",X"FF",X"20",X"0F",X"12",X"7F",X"7F",X"03",X"00",X"00",X"00",X"01",
		X"13",X"00",X"00",X"04",X"1F",X"FF",X"20",X"0F",X"12",X"7F",X"7F",X"01",X"00",X"0A",X"1D",X"12",
		X"23",X"00",X"00",X"FF",X"01",X"FF",X"20",X"0F",X"10",X"88",X"01",X"01",X"00",X"0A",X"1D",X"FC",
		X"23",X"00",X"00",X"FF",X"01",X"FF",X"20",X"0F",X"10",X"92",X"02",X"00",X"01",X"0A",X"0A",X"F3",
		X"08",X"10",X"FB",X"E5",X"31",X"03",X"20",X"0B",X"11",X"78",X"00",X"01",X"00",X"1C",X"12",X"F2",
		X"03",X"E8",X"08",X"0D",X"1C",X"55",X"16",X"15",X"1C",X"4F",X"00",X"01",X"00",X"1C",X"12",X"F2",
		X"0C",X"E8",X"08",X"0D",X"1C",X"55",X"21",X"15",X"1A",X"4B",X"00",X"03",X"00",X"1C",X"12",X"F3",
		X"01",X"E8",X"08",X"0D",X"1C",X"55",X"16",X"15",X"1C",X"32",X"00",X"02",X"00",X"00",X"00",X"E0",
		X"06",X"0C",X"08",X"57",X"01",X"03",X"26",X"F7",X"91",X"1B",X"00",X"EE",X"89",X"EF",X"93",X"ED",
		X"6A",X"00",X"3F",X"EF",X"16",X"EF",X"D5",X"ED",X"0A",X"00",X"1F",X"EE",X"89",X"EF",X"A3",X"ED",
		X"6A",X"00",X"3F",X"EE",X"89",X"F0",X"FB",X"ED",X"4A",X"00",X"1F",X"EE",X"89",X"F1",X"2B",X"ED",
		X"4A",X"00",X"1F",X"EE",X"89",X"F1",X"4B",X"ED",X"4A",X"00",X"1F",X"EE",X"89",X"F2",X"2B",X"ED",
		X"4A",X"00",X"1F",X"EE",X"89",X"F2",X"3B",X"ED",X"4A",X"00",X"1F",X"EE",X"89",X"F0",X"EB",X"ED",
		X"4A",X"00",X"1F",X"EE",X"89",X"F2",X"1B",X"ED",X"4A",X"00",X"1F",X"EE",X"89",X"F1",X"7B",X"ED",
		X"4A",X"00",X"1F",X"EE",X"89",X"F1",X"1B",X"ED",X"4A",X"00",X"1F",X"EE",X"89",X"EF",X"E5",X"ED",
		X"0A",X"00",X"1F",X"EE",X"89",X"F0",X"49",X"ED",X"AA",X"00",X"1F",X"EE",X"89",X"F1",X"5B",X"ED",
		X"4A",X"00",X"1F",X"EE",X"89",X"F1",X"EB",X"ED",X"CA",X"00",X"1F",X"EE",X"89",X"F1",X"FB",X"ED",
		X"CA",X"00",X"1F",X"EE",X"89",X"F2",X"0B",X"ED",X"CA",X"00",X"1F",X"EE",X"89",X"EF",X"5D",X"ED",
		X"0A",X"00",X"1F",X"EE",X"89",X"EF",X"6F",X"ED",X"0A",X"00",X"1F",X"EE",X"89",X"EF",X"81",X"ED",
		X"0A",X"00",X"1F",X"EE",X"89",X"EF",X"B3",X"ED",X"0A",X"00",X"1F",X"EE",X"89",X"EF",X"F5",X"ED",
		X"4A",X"00",X"1F",X"EE",X"89",X"F0",X"9B",X"ED",X"4A",X"00",X"1F",X"EE",X"89",X"F0",X"29",X"ED",
		X"4A",X"00",X"1F",X"EE",X"89",X"F0",X"AB",X"ED",X"4A",X"00",X"1F",X"EE",X"89",X"F0",X"39",X"ED",
		X"4A",X"00",X"1F",X"EE",X"89",X"F1",X"CB",X"ED",X"CA",X"00",X"1F",X"EE",X"89",X"F1",X"DB",X"ED",
		X"CA",X"00",X"1F",X"EF",X"2B",X"F0",X"89",X"ED",X"0A",X"00",X"1F",X"EE",X"8E",X"F0",X"89",X"ED",
		X"0A",X"00",X"1F",X"EE",X"89",X"F0",X"BB",X"ED",X"4A",X"00",X"1F",X"EE",X"89",X"F0",X"CB",X"ED",
		X"4A",X"00",X"1F",X"EE",X"89",X"F0",X"07",X"ED",X"4A",X"00",X"1F",X"EE",X"89",X"F0",X"DB",X"ED",
		X"4A",X"00",X"1F",X"EE",X"89",X"F2",X"4B",X"ED",X"4A",X"00",X"1F",X"EE",X"F5",X"F0",X"79",X"ED",
		X"0A",X"00",X"1F",X"EE",X"89",X"F1",X"3B",X"ED",X"4A",X"00",X"1F",X"EE",X"89",X"F1",X"1B",X"ED",
		X"4A",X"00",X"1F",X"EE",X"89",X"F1",X"6B",X"ED",X"4A",X"00",X"1F",X"EE",X"89",X"F1",X"2B",X"ED",
		X"4A",X"00",X"1F",X"EE",X"89",X"F1",X"4B",X"ED",X"4A",X"00",X"1F",X"EF",X"01",X"F0",X"79",X"ED",
		X"0A",X"00",X"1F",X"EF",X"0D",X"F0",X"79",X"ED",X"0A",X"00",X"1F",X"EE",X"89",X"F1",X"8B",X"ED",
		X"4A",X"00",X"1F",X"EE",X"89",X"F1",X"9B",X"ED",X"4A",X"00",X"1F",X"EE",X"89",X"F1",X"AB",X"ED",
		X"4A",X"00",X"1F",X"EE",X"89",X"F1",X"BB",X"ED",X"4A",X"00",X"1F",X"EE",X"89",X"EF",X"C5",X"ED",
		X"0A",X"00",X"1F",X"EE",X"89",X"F1",X"0B",X"ED",X"4A",X"00",X"1F",X"01",X"09",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"13",X"00",X"FF",X"7F",X"0D",X"1E",X"00",X"00",X"FF",X"00",X"00",X"04",
		X"02",X"10",X"00",X"FF",X"7F",X"0D",X"24",X"00",X"00",X"FF",X"00",X"00",X"04",X"02",X"10",X"00",
		X"FF",X"7F",X"0D",X"32",X"00",X"00",X"FF",X"00",X"00",X"04",X"02",X"10",X"00",X"FF",X"7F",X"0D",
		X"3C",X"00",X"00",X"FF",X"00",X"00",X"04",X"02",X"10",X"00",X"1E",X"00",X"0D",X"76",X"00",X"00",
		X"FF",X"00",X"00",X"04",X"02",X"10",X"00",X"07",X"00",X"04",X"7C",X"08",X"C9",X"FF",X"FE",X"FC",
		X"04",X"02",X"00",X"20",X"1E",X"00",X"0F",X"06",X"02",X"F7",X"09",X"66",X"34",X"01",X"00",X"00",
		X"00",X"F9",X"42",X"0F",X"06",X"02",X"F7",X"09",X"DF",X"D9",X"01",X"00",X"00",X"00",X"F9",X"42",
		X"14",X"08",X"02",X"F7",X"FF",X"DF",X"D9",X"00",X"00",X"00",X"00",X"FF",X"8F",X"15",X"08",X"02",
		X"F7",X"FF",X"DF",X"D9",X"00",X"00",X"10",X"00",X"FF",X"8F",X"F4",X"6D",X"14",X"09",X"02",X"F7",
		X"FF",X"DF",X"D9",X"00",X"00",X"10",X"00",X"FF",X"8F",X"F4",X"8B",X"14",X"0A",X"02",X"F7",X"FF",
		X"DF",X"D9",X"00",X"00",X"10",X"00",X"FF",X"8F",X"F4",X"9A",X"14",X"08",X"02",X"F7",X"FF",X"DF",
		X"D9",X"00",X"00",X"10",X"00",X"FF",X"8F",X"F4",X"6D",X"08",X"08",X"02",X"F7",X"FF",X"DF",X"D9",
		X"00",X"00",X"00",X"00",X"80",X"04",X"14",X"09",X"02",X"F7",X"FF",X"DF",X"D9",X"00",X"00",X"00",
		X"00",X"FD",X"8F",X"F4",X"C5",X"14",X"0A",X"02",X"F7",X"FF",X"DF",X"D9",X"00",X"00",X"00",X"00",
		X"F8",X"88",X"F4",X"D4",X"14",X"09",X"02",X"F7",X"FF",X"DF",X"D9",X"00",X"00",X"00",X"00",X"FD",
		X"88",X"F4",X"E3",X"14",X"08",X"02",X"F7",X"FF",X"DF",X"D9",X"00",X"00",X"00",X"00",X"FF",X"8A",
		X"F4",X"A9",X"01",X"02",X"04",X"FF",X"40",X"FF",X"3F",X"00",X"00",X"10",X"00",X"FF",X"FF",X"F4",
		X"F2",X"01",X"02",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",X"10",X"00",X"FF",X"FF",X"F5",X"01",
		X"01",X"04",X"00",X"00",X"00",X"FF",X"00",X"01",X"03",X"11",X"00",X"FF",X"FF",X"F5",X"10",X"08",
		X"13",X"02",X"F9",X"FF",X"E3",X"E0",X"05",X"08",X"14",X"00",X"C0",X"05",X"01",X"00",X"01",X"01",
		X"FF",X"D9",X"55",X"00",X"00",X"10",X"00",X"00",X"00",X"01",X"00",X"01",X"01",X"FF",X"D9",X"55",
		X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"00",X"01",X"01",X"FF",X"D9",X"55",X"00",X"00",X"12",
		X"00",X"00",X"00",X"01",X"00",X"01",X"01",X"FF",X"D9",X"55",X"00",X"00",X"13",X"00",X"00",X"00",
		X"01",X"00",X"01",X"01",X"FF",X"D9",X"55",X"00",X"00",X"14",X"00",X"00",X"00",X"02",X"06",X"04",
		X"02",X"FF",X"00",X"00",X"00",X"00",X"10",X"00",X"FF",X"7F",X"37",X"01",X"00",X"00",X"FF",X"00",
		X"00",X"02",X"01",X"11",X"00",X"FF",X"7F",X"0A",X"05",X"00",X"09",X"FF",X"83",X"DE",X"00",X"00",
		X"10",X"00",X"FF",X"FF",X"F5",X"87",X"01",X"04",X"02",X"13",X"FF",X"1E",X"63",X"00",X"00",X"10",
		X"00",X"FF",X"03",X"F0",X"05",X"02",X"16",X"FF",X"82",X"94",X"00",X"00",X"10",X"00",X"FF",X"7F",
		X"02",X"0F",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"02",X"18",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"04",X"14",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"FB",X"00",X"01",X"07",X"06",X"DF",X"F2",X"05",X"03",
		X"14",X"00",X"FF",X"00",X"F5",X"E6",X"FB",X"00",X"01",X"07",X"06",X"DF",X"F2",X"05",X"03",X"14",
		X"01",X"FF",X"00",X"F5",X"F5",X"FB",X"00",X"01",X"07",X"06",X"DF",X"F2",X"05",X"03",X"14",X"02",
		X"FF",X"00",X"F6",X"04",X"FB",X"00",X"01",X"07",X"06",X"DF",X"F2",X"05",X"03",X"14",X"03",X"FF",
		X"00",X"F6",X"13",X"FB",X"00",X"01",X"07",X"06",X"DF",X"F2",X"05",X"03",X"14",X"04",X"FF",X"00",
		X"F5",X"D7",X"01",X"02",X"01",X"01",X"FF",X"D9",X"55",X"F7",X"01",X"11",X"00",X"FF",X"7F",X"21",
		X"02",X"FF",X"0E",X"00",X"01",X"01",X"00",X"C7",X"11",X"00",X"FF",X"7F",X"21",X"02",X"FF",X"0E",
		X"00",X"01",X"01",X"00",X"D3",X"11",X"00",X"93",X"80",X"F6",X"4B",X"4A",X"03",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"11",X"00",X"0F",X"80",X"F6",X"4B",X"02",X"02",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"15",X"11",X"00",X"FF",X"7F",X"04",X"01",X"00",X"00",X"FF",X"00",X"00",X"01",X"01",
		X"11",X"00",X"FF",X"7F",X"01",X"01",X"00",X"00",X"FF",X"00",X"00",X"00",X"E3",X"11",X"00",X"FF",
		X"7F",X"01",X"06",X"00",X"00",X"FF",X"00",X"00",X"01",X"35",X"11",X"00",X"FF",X"7F",X"01",X"0B",
		X"00",X"02",X"00",X"00",X"00",X"01",X"FA",X"01",X"00",X"FF",X"7F",X"01",X"0B",X"00",X"02",X"FF",
		X"00",X"00",X"01",X"ED",X"11",X"00",X"FF",X"7F",X"01",X"0B",X"00",X"02",X"FF",X"00",X"00",X"01",
		X"EB",X"11",X"00",X"FF",X"7F",X"01",X"0B",X"00",X"02",X"FF",X"00",X"00",X"01",X"DE",X"11",X"00",
		X"FF",X"7F",X"01",X"0B",X"00",X"02",X"FF",X"00",X"00",X"01",X"C7",X"11",X"00",X"FF",X"7F",X"01",
		X"0B",X"00",X"02",X"00",X"00",X"00",X"00",X"F0",X"11",X"00",X"40",X"00",X"01",X"0B",X"01",X"03",
		X"01",X"01",X"02",X"01",X"EE",X"11",X"00",X"40",X"00",X"3C",X"02",X"01",X"03",X"01",X"01",X"02",
		X"01",X"FF",X"12",X"DD",X"40",X"00",X"01",X"0B",X"01",X"03",X"01",X"01",X"02",X"01",X"EE",X"11",
		X"00",X"10",X"80",X"F7",X"05",X"01",X"0B",X"00",X"02",X"00",X"00",X"00",X"00",X"F0",X"11",X"00",
		X"40",X"00",X"01",X"0B",X"01",X"03",X"01",X"01",X"02",X"01",X"EE",X"11",X"00",X"10",X"80",X"F7",
		X"21",X"01",X"0B",X"00",X"02",X"FF",X"00",X"00",X"01",X"C7",X"11",X"00",X"FF",X"7F",X"07",X"04",
		X"00",X"02",X"00",X"04",X"07",X"7F",X"FF",X"13",X"01",X"13",X"00",X"FF",X"7F",X"0C",X"02",X"01",
		X"0B",X"FF",X"00",X"00",X"00",X"BE",X"11",X"00",X"FF",X"7F",X"0C",X"05",X"01",X"0B",X"FF",X"00",
		X"00",X"00",X"BE",X"01",X"00",X"FF",X"7F",X"08",X"02",X"00",X"00",X"D4",X"00",X"00",X"01",X"EF",
		X"11",X"00",X"81",X"00",X"02",X"01",X"00",X"01",X"D7",X"01",X"01",X"01",X"F4",X"13",X"03",X"2D",
		X"00",X"01",X"09",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"03",X"00",X"FF",X"00",X"02",X"01",
		X"00",X"00",X"20",X"00",X"00",X"00",X"35",X"01",X"00",X"81",X"01",X"01",X"02",X"05",X"00",X"FF",
		X"00",X"00",X"F9",X"FA",X"11",X"00",X"FF",X"FF",X"F7",X"9A",X"02",X"02",X"00",X"00",X"FF",X"00",
		X"00",X"46",X"7D",X"11",X"00",X"FF",X"FF",X"F7",X"8B",X"03",X"74",X"02",X"04",X"04",X"DC",X"DB",
		X"FB",X"08",X"14",X"FB",X"FF",X"0F",X"03",X"74",X"02",X"04",X"04",X"DC",X"DB",X"FB",X"08",X"14",
		X"F8",X"FF",X"0F",X"03",X"74",X"02",X"04",X"04",X"DC",X"DB",X"FB",X"08",X"14",X"F9",X"FF",X"0F",
		X"03",X"74",X"02",X"04",X"04",X"DC",X"DB",X"FB",X"08",X"14",X"FA",X"FF",X"0F",X"03",X"74",X"02",
		X"04",X"04",X"DC",X"DB",X"FB",X"08",X"14",X"02",X"FF",X"0F",X"09",X"05",X"08",X"F7",X"FF",X"DF",
		X"D9",X"00",X"02",X"00",X"00",X"80",X"04",X"09",X"05",X"09",X"F7",X"FF",X"DF",X"D9",X"00",X"02",
		X"00",X"00",X"80",X"04",X"09",X"05",X"0A",X"F7",X"FF",X"DF",X"D9",X"00",X"02",X"00",X"00",X"80",
		X"04",X"0A",X"02",X"01",X"0B",X"FF",X"00",X"00",X"00",X"BE",X"12",X"00",X"FF",X"7F",X"0A",X"02",
		X"07",X"0E",X"05",X"03",X"03",X"03",X"C3",X"10",X"00",X"FF",X"03",X"04",X"3B",X"00",X"00",X"FF",
		X"00",X"00",X"04",X"02",X"10",X"00",X"FF",X"7F",X"06",X"4C",X"00",X"00",X"FF",X"00",X"00",X"04",
		X"02",X"10",X"00",X"12",X"00",X"06",X"86",X"00",X"00",X"FF",X"00",X"00",X"04",X"02",X"10",X"00",
		X"08",X"00",X"06",X"26",X"00",X"00",X"FF",X"00",X"00",X"04",X"02",X"10",X"00",X"0A",X"00",X"06",
		X"1F",X"00",X"00",X"FF",X"00",X"00",X"04",X"02",X"10",X"00",X"08",X"00",X"06",X"1E",X"00",X"00",
		X"FF",X"00",X"00",X"04",X"02",X"10",X"00",X"FF",X"7F",X"06",X"1D",X"00",X"00",X"FF",X"00",X"00",
		X"04",X"02",X"10",X"00",X"2F",X"00",X"08",X"19",X"00",X"00",X"FF",X"00",X"00",X"04",X"02",X"10",
		X"00",X"08",X"00",X"21",X"02",X"FF",X"0E",X"00",X"01",X"01",X"00",X"D3",X"11",X"00",X"FF",X"8F",
		X"F8",X"A2",X"01",X"0B",X"00",X"02",X"00",X"00",X"00",X"00",X"F0",X"11",X"00",X"40",X"80",X"F8",
		X"B1",X"21",X"02",X"FF",X"0E",X"00",X"01",X"01",X"00",X"D3",X"11",X"00",X"FF",X"7F",X"0D",X"1E",
		X"00",X"00",X"FF",X"00",X"00",X"04",X"02",X"10",X"00",X"0C",X"00",X"0D",X"24",X"00",X"00",X"FF",
		X"00",X"00",X"04",X"02",X"10",X"00",X"FF",X"7F",X"0D",X"32",X"00",X"00",X"FF",X"00",X"00",X"04",
		X"02",X"10",X"00",X"FF",X"7F",X"0D",X"3C",X"00",X"00",X"FF",X"00",X"00",X"04",X"02",X"10",X"00",
		X"FF",X"7F",X"04",X"3B",X"00",X"00",X"FF",X"00",X"00",X"04",X"02",X"10",X"00",X"FF",X"7F",X"06",
		X"1C",X"00",X"00",X"FF",X"00",X"00",X"04",X"02",X"10",X"00",X"19",X"00",X"09",X"24",X"00",X"00",
		X"01",X"E3",X"F5",X"04",X"02",X"10",X"00",X"11",X"00",X"09",X"24",X"00",X"00",X"01",X"E3",X"0E",
		X"04",X"02",X"10",X"00",X"0D",X"00",X"0B",X"32",X"00",X"00",X"FF",X"6A",X"0F",X"06",X"02",X"10",
		X"00",X"FF",X"7F",X"04",X"3B",X"00",X"00",X"FF",X"00",X"00",X"04",X"02",X"10",X"00",X"43",X"00",
		X"04",X"3B",X"00",X"00",X"FF",X"00",X"00",X"04",X"02",X"10",X"00",X"33",X"00",X"04",X"3B",X"00",
		X"00",X"FF",X"00",X"00",X"04",X"02",X"10",X"00",X"08",X"00",X"04",X"3B",X"00",X"00",X"FF",X"00",
		X"00",X"04",X"02",X"10",X"00",X"33",X"80",X"F9",X"4D",X"09",X"23",X"00",X"00",X"01",X"E3",X"0E",
		X"06",X"04",X"10",X"00",X"0D",X"00",X"08",X"26",X"00",X"00",X"01",X"E3",X"0E",X"06",X"04",X"10",
		X"00",X"0D",X"00",X"08",X"26",X"00",X"00",X"01",X"E3",X"0E",X"06",X"04",X"30",X"00",X"0D",X"00",
		X"06",X"1C",X"00",X"00",X"FF",X"00",X"00",X"04",X"02",X"30",X"00",X"19",X"00",X"09",X"24",X"00",
		X"00",X"01",X"E3",X"F5",X"04",X"02",X"30",X"00",X"11",X"00",X"09",X"24",X"00",X"00",X"01",X"E3",
		X"0E",X"04",X"02",X"30",X"00",X"0D",X"00",X"EE",X"28",X"F4",X"60",X"ED",X"EE",X"F6",X"4B",X"ED",
		X"EE",X"F7",X"57",X"ED",X"EE",X"F7",X"64",X"ED",X"EE",X"F7",X"9A",X"EE",X"54",X"F7",X"4A",X"EE",
		X"12",X"F4",X"6D",X"EE",X"3C",X"F4",X"A9",X"EE",X"00",X"F5",X"10",X"ED",X"EE",X"F7",X"3D",X"ED",
		X"EE",X"F6",X"5A",X"ED",X"EE",X"F6",X"74",X"ED",X"EE",X"F6",X"81",X"EE",X"34",X"F6",X"8E",X"ED",
		X"EE",X"F6",X"CF",X"ED",X"EE",X"F6",X"DC",X"ED",X"EE",X"F6",X"E9",X"ED",X"EE",X"F6",X"2F",X"ED",
		X"EE",X"F6",X"3C",X"ED",X"EE",X"F3",X"EB",X"ED",X"EE",X"F3",X"F8",X"ED",X"EE",X"F4",X"05",X"ED",
		X"EE",X"F4",X"12",X"ED",X"EE",X"F4",X"1F",X"ED",X"EE",X"F4",X"2C",X"ED",X"F2",X"F4",X"39",X"ED",
		X"F8",X"F4",X"39",X"ED",X"EE",X"F7",X"8B",X"ED",X"EE",X"F6",X"67",X"EE",X"48",X"F6",X"67",X"EE",
		X"62",X"F7",X"4A",X"EE",X"12",X"F5",X"1F",X"EE",X"00",X"F5",X"6D",X"ED",X"EE",X"F5",X"87",X"EE",
		X"12",X"F4",X"A9",X"ED",X"EE",X"F6",X"9B",X"ED",X"EE",X"F6",X"A8",X"ED",X"EE",X"F6",X"C2",X"ED",
		X"EE",X"F6",X"F6",X"ED",X"EE",X"F7",X"12",X"ED",X"EE",X"F7",X"A9",X"ED",X"EE",X"F7",X"B6",X"ED",
		X"EE",X"F7",X"C3",X"ED",X"EE",X"F7",X"D0",X"ED",X"EE",X"F7",X"DD",X"ED",X"EE",X"F7",X"EA",X"ED",
		X"EE",X"F7",X"F7",X"ED",X"EE",X"F8",X"04",X"ED",X"EE",X"F8",X"11",X"ED",X"EE",X"F8",X"1E",X"ED",
		X"EE",X"F8",X"2B",X"ED",X"EE",X"F8",X"38",X"ED",X"EE",X"F8",X"45",X"ED",X"EE",X"F8",X"52",X"ED",
		X"EE",X"F8",X"5F",X"ED",X"EE",X"F8",X"6C",X"ED",X"EE",X"F8",X"79",X"ED",X"EE",X"F8",X"86",X"ED",
		X"EE",X"F8",X"93",X"ED",X"EE",X"F8",X"BE",X"ED",X"EE",X"F8",X"CB",X"ED",X"EE",X"F8",X"D8",X"ED",
		X"EE",X"F8",X"E5",X"ED",X"EE",X"F8",X"F2",X"ED",X"EE",X"F8",X"FF",X"ED",X"EE",X"F9",X"0C",X"ED",
		X"EE",X"F9",X"19",X"ED",X"EE",X"F9",X"26",X"ED",X"EE",X"F9",X"33",X"ED",X"EE",X"F9",X"40",X"ED",
		X"EE",X"F9",X"4D",X"ED",X"EE",X"F9",X"5A",X"ED",X"EE",X"F9",X"69",X"ED",X"EE",X"F9",X"76",X"ED",
		X"EE",X"F9",X"83",X"ED",X"EE",X"F9",X"90",X"ED",X"EE",X"F9",X"9D",X"ED",X"EE",X"F9",X"AA",X"1C",
		X"80",X"40",X"29",X"1B",X"10",X"09",X"06",X"04",X"07",X"0C",X"12",X"1E",X"30",X"49",X"A4",X"C9",
		X"DF",X"EB",X"F6",X"FB",X"FF",X"FF",X"FB",X"F5",X"EA",X"DD",X"C7",X"9B",X"10",X"00",X"F4",X"00",
		X"E8",X"00",X"DC",X"00",X"E2",X"00",X"DC",X"00",X"E8",X"00",X"F4",X"00",X"00",X"20",X"4C",X"45",
		X"41",X"41",X"43",X"47",X"77",X"87",X"90",X"97",X"A1",X"A7",X"AE",X"B5",X"B8",X"BC",X"BE",X"BF",
		X"C1",X"C2",X"C2",X"C2",X"C1",X"BF",X"BE",X"BB",X"B6",X"B1",X"AC",X"A4",X"9E",X"93",X"10",X"3C",
		X"10",X"17",X"3F",X"70",X"92",X"95",X"7F",X"7C",X"7E",X"8A",X"BE",X"E7",X"EF",X"C5",X"7F",X"08",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"10",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"48",X"8A",X"95",X"A0",X"AB",X"B5",X"BF",
		X"C8",X"D1",X"DA",X"E1",X"E8",X"EE",X"F3",X"F7",X"FB",X"FD",X"FE",X"FF",X"FE",X"FD",X"FB",X"F7",
		X"F3",X"EE",X"E8",X"E1",X"DA",X"D1",X"C8",X"BF",X"B5",X"AB",X"A0",X"95",X"8A",X"7F",X"75",X"6A",
		X"5F",X"54",X"4A",X"40",X"37",X"2E",X"25",X"1E",X"17",X"11",X"0C",X"08",X"04",X"02",X"01",X"00",
		X"01",X"02",X"04",X"08",X"0C",X"11",X"17",X"1E",X"25",X"2E",X"37",X"40",X"4A",X"54",X"5F",X"6A",
		X"75",X"7F",X"73",X"20",X"00",X"00",X"00",X"04",X"00",X"A3",X"11",X"00",X"01",X"01",X"10",X"04",
		X"FF",X"12",X"14",X"01",X"01",X"04",X"14",X"3D",X"53",X"01",X"01",X"01",X"02",X"18",X"01",X"14",
		X"00",X"00",X"00",X"08",X"1A",X"81",X"25",X"00",X"00",X"00",X"16",X"22",X"01",X"16",X"01",X"01",
		X"01",X"01",X"38",X"FE",X"10",X"00",X"00",X"00",X"20",X"4C",X"F1",X"10",X"00",X"00",X"00",X"4D",
		X"4C",X"F1",X"15",X"00",X"00",X"00",X"4D",X"4C",X"F1",X"16",X"00",X"00",X"00",X"4D",X"4C",X"FE",
		X"10",X"00",X"00",X"00",X"20",X"4C",X"08",X"10",X"20",X"30",X"14",X"18",X"20",X"30",X"40",X"50",
		X"40",X"30",X"20",X"10",X"0C",X"0A",X"08",X"07",X"06",X"05",X"01",X"02",X"02",X"03",X"98",X"90",
		X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"01",X"01",X"02",X"02",X"04",X"04",X"08",X"08",
		X"10",X"20",X"28",X"30",X"38",X"40",X"48",X"50",X"60",X"70",X"80",X"A0",X"B0",X"C0",X"08",X"40",
		X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",
		X"08",X"40",X"01",X"01",X"01",X"02",X"02",X"03",X"03",X"04",X"02",X"02",X"03",X"03",X"04",X"04",
		X"05",X"03",X"03",X"03",X"04",X"04",X"05",X"05",X"06",X"02",X"02",X"02",X"03",X"03",X"04",X"04",
		X"05",X"03",X"03",X"03",X"04",X"04",X"05",X"05",X"06",X"04",X"04",X"04",X"05",X"05",X"06",X"06",
		X"07",X"07",X"07",X"07",X"08",X"08",X"09",X"09",X"0A",X"0C",X"0C",X"0C",X"0D",X"0D",X"0E",X"0E",
		X"0F",X"06",X"06",X"06",X"07",X"07",X"08",X"08",X"09",X"02",X"02",X"02",X"03",X"03",X"04",X"04",
		X"05",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E9",X"B9",X"E0",X"01",X"E9",X"DD",X"E0",X"01");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
